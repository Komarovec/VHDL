`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m+Mk59EAMaEvcL8Kwbptjru+lm/NMyOFpKdEsAYieekU9TohoTFJSeX4Qy0MCm3bSmSfFaijpNrx
pCdds3c7Mw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eaV6HPOXe9nLJXggg6KOmcxYvFLPnlZVlD2veVPfuEDrvqcpIeflxbrtfilnOYqpg1R+tAKtClqE
pvzxfboR06Mp+ULbBkBvVkB7b4pgDBGUlECQJB+oE8vVv6Ord9+iXdoqBiVyg+GbkVzqHaxsN7O/
icKe2PWre0gvWhz0yvU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AsNm91ZG4N2uiVr32mJCQ31e7MRRPElAnC4WlDK8TXPTud+OpVlnpwiJaEfGQZnQp3mkFmZlbFpV
D/XKy9J7eeGBrJ3m7JU0EV43CzzpPyBWK8+mUqVoX/vUCh/G02OpOoNkXBU8XMCkZSy2OKzHliVR
QVwDpxfi1hyu54IzzwI/t73POzXIMrVoDVaRxAPSFIOWJGjqkBgjhr9fv98FysH0qEnWbIRGjoQm
2+exctbpfPZ7UPQhAjXT9dOidD9FGOAJ56g3vk8xgrXandychs3NlIr+mC3ZjqcBjKagN3IULEhg
N+5EIRHqyFPHYuvFPnNUq7YnA2NSZrYqtLndjQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KUl60kFJoHCucCRs5dtQAH6iwMTh9jKT09SW6/cFFfp8nQubb3fiBfJU9gYSrSbNxO5ElkGZMvT6
f3xU1dlUzmSdP2cm5SSjnKg4MzI2q7kDm2hQ7i38PTGMX+JOekIwd2nuf8ik/Ugg9VEe++sFOq3E
G3PBBL1bzbOwoqNYMKXfyKDTVwGU2Ug15246OIDB98wnIBIUDygszsQqSRe9F8pbjfHm2QL0hu15
AYPDcthUfnAOdTqDh6MGuaSR1NNPoMCYXECihWSfAy96mgFMxnDLXAxjv66NxPMchhcW8oZHD/r4
MZv9qj7k85mHLS64sFtdqgdSsNToqPXhwF8R9Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iHD41KTQE10umuJdb95an5zAG3dQOcP4qYjzX6HT865+ghStilUvaQMQGndrQVlfAP/yAdoHTwO4
9VCl26hube7oz0QCgG1a0KxRYEUXkdvnv/xQt1Mojeyg0Uc9EOd5/OFkiQwMu42cl2nejxYllMIC
1UyCrrVetqTCZLb+XQ0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RAdeOZjyJxieb6py2nKEFYXKyKy6WrDcHlFQBf6f08MWEzyWpXcOY4jBxDXORRI8OaaNerjVHRDY
Auj3duVBWPw5GWqT7r/pbieD4FkzLNpANF9DMnQhTxMcAwiiNp5fzFxJucMVgPAj4iB6GS8NBejn
7lmS9x72ZHk7zIP0Yej4vqmdy76XldyoDCdR3RET4UsXYOjbhr4qvkq0RHHNQry1BEzWwtQ67hTX
IkObOUf+nGKWF6E9LWCBvqBi2aHtt+4RVuQ4tVQvczyjkmrjD0iLeZEg5suY98kF0iquwJGJhXmB
jXPjY89FANu+is4sEK/lzUa32QDcTksQkEkTqQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WfZnhPbtwOwgBWtxF6/ewwvNGTS+NBvjGA9tsxe8SIeHv3Y+kMzquM1CwwcmPKk7ljPPK8k/UULb
pkGd8d/M2NUlLc3ULMQi4NZZEuu/lRndWXp3/KLqxx9/Sb3yuq7F0pRB59Yv3HdHS3tkLnAnjY+f
GgKPOC3Mx2teEQ4NSNRYBFJbKwP8dd5/a7WcqBxGXSh7bsfECLRuAOkgYEa5B6Xo3Q6ZWk1tLPgG
sN8Py0/f/ULiaUGwvmLfSzlUCjCjkjXsQrz60L87tnQ4gGkfMreGgJC66ZKYMUNKlTdlBdL7TMrB
KNo/NXwB8ws6eqNTvo55GPKDdEBuD6do26wFdA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
siwW7+1Pu/HvZtOOT8oIJ2sQIaFE8o53vAuBib7YwKonCOiopn1iFJiZSmUK+Sz2KTaD5UxDjBwe
OHSH/dQW1eLH229I2dFK1LSzKn8ccuQNaiZ17dE0JIWKagXClEuQDDrlQICj90ov9XOHSgUYV+bi
wTp1qa02gULZ96jPjRE3rFC5PHPExCZPDI45cef+4KxXMBLDktr6+ll/VH4g2JBmBAxfjLEQED7b
lsw3hrlxYS1mWpcSHp47pfkjyibK2fGrrV/+oSA4fTbhROBQaUfwW4vp2wxHuuu1WR6mzNaTvHuO
qd0Nnvv42i1iVQz5naiY5p4BHQnH+1aFA0fI6Q==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XQlnW7KBXb5ghdFrIj3e+hc0/c9PA/o3Ztn5NJ3YC5+EKeWROXnw9dD4P+CTnl7W/o6wjCO/ImwM
r6kLgua2sNFHO/72vUzwLtl+RwPLgYbHisZlxwnIOhuWqqqQla0UgsO+lrjZd/llIF5mGABk2xzi
lObHqIiHva3ry4rc1NOwo03xbvsJKdgTAxeWmJCy/Y7pt4rpWFE1fQzkPgIPoX6R+jLlr5EtMbyW
JEhdmPYlKZjdjVeSDcZMREIYNNGiaPv+T4OjaWUGXQOcgK0uZ1FdHufgjX7LrMP4xLtaWeoi1skv
ttlWhLx6q8DF/7Fmli75scOIJHmAaH/Q66zpww==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 183840)
`protect data_block
ec4qH+rSlyFgSEY1SJhIOVhXda5tlG2Qp1litayxn696aSc9uU0dGTDskaZR9RZByWEZebPGGZPu
+bGwwehKsQQp8JsRfuSxJIoVxib5sluN5hgoPVNxIbv9Z23EACDA++GqGP6kyH/Z4Dih+fpV+Iv6
08eppOMh9v5rcohC5IHljaRCUcgSykiNHyh/m+DqiCF08FWYd8v6zaunkxE08bfLjG/VETb0bzog
ViV2OEagRTlAiJH85Lae/ttFN860C1NqmKCqppY8vpjbNDezsecR3R6Qct68x6wrP8s2weA9v/Hw
jeCL6ShbzHiYoqowGkL1L6OpLBCo0lj9lJayoUaHqZIMDtJ68dctjckSoNIHteScwCR9JsR7nCon
sBBIzwyJQowRoZvhJ/Bsid171fo0Ik8IG6+zIwg4BV/rvb3qTmAp7tXkc2Xbtmau+5xgJTMX/iHJ
Z5y18yUsW7rx21wUWAd76B7n8izBVGqVuC+mF6CBUJBgvZ7aeTDmDnpPksyn5yGQ4H6HAl8dswJC
AswOVKm0VflWDcgiE8K3ubmMWnA+EoZ/AL4UdAbIp5i3ZOrvjf+H3x7QpMgR2l1m9Cmj92JoVEwH
i7rwgxenQOLEayauw7ruR4TR52LMNl11qZ2Ya2humJfNsni2zSoB5CYAScQugPgWF02ImvbfRcmh
6R3SrOGRSGLKzrhv4EF5td9WqDYXBJEDf8Oe0H9r3XJ5w3gRdHNYd44pUGmIc2EQdraoIh6YkBC+
73sVfJu/mG6pTVF+gotEU8gfZ+fMWgxWFV5MZlF9r4rRkx4EwVbq5TdJDhBd6WTRnu6ardEET/aD
sLuwHEMLc5yZtmcKQULonCGcC3OL+3GOi+CN4sVV3boNZMB6IQYNubVDX0e3z27bdW9FJb8kYZJ7
uI7gqgp6DmopIKJaVM9Gg7NQUrQTvGCESF2adamWk7xpRvnbJxVicRJ7q+mojDaxYxmogQaRCUGb
lEkzeaeodEWIeWleildCyrNkPF9g+26AEmFhXdj/kzudAVRt2TXslP6sle8K+hhdf9NTSzNlD5xf
lRkT9UDVH+Wpb0PgEogsNPSro3zLSmIlh3Sb0nbcTdIpuw5a+AH89727b2EmwpJs3PtUIknFOz4I
Vm983TviIiQkgmuQ9zCZ3O2Eox1SgiKy7IHsTNUFSM4Inr/zJuUTHZFyIEACWyFqskMQinQS60yY
eytxu9Gr6cZiEFFVZPwqVMJsqbmPgTB0Zurb2ZaeFyA7nnKCQVPgeRLoWuNmdsjJ73gJXDgBvLHo
3WykqQNIQx4E4HiahjqSB4ITXLnyTinJ87e0vFGbpqlNEG6geLB3+s3/aDmkEQFRaGtDahk8Pl5p
tDkpCr3252QtvjPGBEy9cjBTBAtKO8aEOHe6ppPCIwTyfO0IgCrJVxOliDSOp8U+d339NIQPZviC
kJvhSviCiMEFgYoOG/GPDQjpUZ+OAN9feCpfeRjOT0gx6zQzgS7V4wuBOyBfNMTZip4MubMDDNpJ
aXR/YjJMIvzRo7NM+z9qkAeW3k24oPlBF19DtxZmNdWQgdBQ76vbhMn0nrKhsy49Fz+g4SG+RZOg
nR6fJ9TgNE2nuA6Zs6iyUuJUKFoaHf1jprMEeeGyYET6N+Pc+V543N58wBjkDHvrPHEyjPYo13zE
0ODTuRVKHrfie88MB7UBt6w12MXrPo9B+YRo6bqSCP+QRnNgoW4nZiWjp+O9ZBIzMp/+aH2VUQst
s+QNuCYDLtirj4U0lCpDoFRLZBKnYmGDv4vfCQfpg4mqTeJmaJeztdEcUqcDKiPNaI+F+R+aRHjo
Dy472Uy0NktWBROj2MJ5ADIPS4uoIoTTtUXfb3U4ygfnZuEDd7akM2sQB9K1ViPTBh5dOz1nHI+3
f39UV19hpo8N2NPbEF9fbzycfZAK00UQTmgdVnm6AREZkshtSU5VW6aH++FLDpkoRA6aNnVL+39x
sI5KqRzfDpO7+v/IsfjciYhji6hhpHEuJwo3AEMyev7oeTWlta5IHV8zjuBXloqsEW59zqJW2hje
XWre2oAu5zxF7fjs9D5DboE72/Pf2D5xdz/ZuTTHnvzzH790YNwwWViIZeVJdqK+lkSCdZCQaTMD
IDshXsKIvKO43CN+zuXOmhLQmtL1iloIjk2hvKHgUWH2m0fEHtRYBiaVRfZpHiAueF6LOEY00TOY
fZYLZ4hQnB4woN9O+RXbkKU5+MxG3T3Ha6dcDVq4mPh8XdxQCCy7vbsFe1IjWjACb8+qlpq++Fh2
YgWglGlI9hRm1Z2Oy0u26ipE6132HVlJxEVl0KrCYwLfFtAVjBQiBtfkyRAdi6WzBcvVCK7Ew+3a
uiFyxn4QRH+gGmOgiaWDBmWlgwn6/9kqNdwbweT9kRueHXx0A6wTLr3zbcISTGCauWqaab0NiUYS
Qxcx6epEm/0ArWEMnPRcOd8/htkWEpgG/h/mqjm+HSUD28H4cUyQ7oWlr+zxHuZY0nIklV2nGDJr
6hu/zMcO2B7lgwsP3wDvfe1P1KZKjYaV/E2IchbEmQQgumMqnoKcL0o39fG9Qmn3N5jX2ldCR0fh
vGl52Lk/BpPw9yE7LyoaMIbWAmJgruOKGIQw/5aiTbGmoPrNxUEFyXEQGCc0wZxyAHxQ0YHThPvz
sSx3uJxGHhu7V0DmT9W8/BKhP5+VZKdG1X1m7JwaHE3pZ3DgeJsC7eK4bCwDPs8ye2+6419AFWUM
wWOD0tUw0XWbQVbcVVQ3FnJSkpgRM2bxlvpgPinujYfnRsupWVrA0MyfkID5arOe2LOMgNsWCbNn
BNPK8Q80CTaYM+D1BbF7uXqzI2qB8TnTh9S+AamFeo/nM/lzjzj632MDaPiWtzLFam+uttySkKNV
09gipsU3P90kauwN3DLHvqHb7yMKzNbBtdRtNi4LAI+Tj1xEPUvR3ZzmcmlMvYoW8VuHcWJYFGKS
6ehP+Jn8NE+J/TtPiGOEB926AsSn+D3UySnea39sVHKh58xIyETuznrw73qy8hiwtrYQhPu3SkNv
htOy1rTEJy6zaqM10hSc72P+zKAae6ye8q3sUzliFpHk9seu31NKjaL23gh5wZc4GrYicbeef82x
8gR7vVnSL+5KQ78Kzx73hJsmB6RMgxhk3CbgfedypFJro6V0ZlX44NPvsWFIBmwPwVdMFtyjA/49
slDhJa/oJ4yNuvpvo59qxgQhm4cJoER2GIZJGlEWtLJFB2fKBO+3QPypRKj/CnbBxn+Y26qVYK6a
uFPuZ83p1PjX5Dpvw8HTKvJu5AnEvCY+iwCwg75QKPRaAumRkVTR70ojEwLXIc3c2ijNg8ED5d9s
+oW0ZLmwHGX02QQarnhBMD8za75FDz6+yvWR+AnJcEp/XI21DUlGSSRHwCdoWo7ZRVMpHXCUDOdc
dzaAFsEHAZSAekbXqvpi+4XYCq7ei9ldWanJLLbP88kLZbojk1i7fyfgd6mFxZei9sQIrXfVO5SP
pYD3MM8BpbYmb81jxgI0ifyU7GGG4w8TmrV8iMsQsX02DwsnOB43TejRengM7Ld741lbGQEe/DP5
J73L67YVgthphWt4eaLDC4lsVMOOwUu1P15cyWP3xLuM2r+lRELX/WIl8ESabtESHSxU958n5xqV
Y8+8cqT3WlN+yHn52v2tZjp26sN9lW8W5xhvzaMuhpZcTULWN8mm0yygKmb7aXHwydQg/VQEAwHk
VN/VRzxd6YER9fEHW1Wtj4zmObJcBdKhIDWVMEMvGqUVA++jNR6qzehB8dMWrGQ/sMrDxxjUxiGe
TjcJB4ZghEeaXAKabMOuqMKaBz062vKnxXZ+kN8c8C1u1NxONI0DtaNLroLsusn/6cpvYE9z55qc
9hkRpsGfEGs+7YSamTaqOoy7Fd8LlcrNObP6s9V5625PSwsrLV8VuaM+Ts3IzJ8jJmFZFqpNU5W8
qbTvpyGPCRrdDUI9D8onWL7jGmkbuDq2Zwc0NgNWsHvZ2o8JxjoVkyFhOJC8LZ4rMsFhHNqy584Y
DkS5tdpQZ9wEUhlqcC690VDWlYX+uTfFyeQwUSg965nXjLeRwmzemuD0GpVxoy37WOBUgll1KmRv
zKoG5krdvEcpYav4yl6uImDPCFeON5eN21msWnI7Y9xAjURfzfziFVRpoFNDlHCIU6hO+uOAaKpY
bae//kmdYln7AXTiaJPhO2eqOhFfh39ifYE9SWH8Yxij0Sb+Xc/juyLdhBvV65uRUR6qLgzxtvxl
XlkVQL6fKhus57Gn3xIUKrQwoVY37YBO5kHe6TykOVRw1ak3mvATsB2P0lOlEV+8ceVgeK/j9FOR
rDntWuFKjsWaN0+Q56/9Bfs4Mf+Iel4DMh3G/jd8uqaI8mAN4TOeYKMBpZsVDfHdCYH2dDYs4ftY
Sz7MRf18vB8aFkiZ+ovyAGB7d8z42v3roktEAVgYiA6rg76YZRi2ju3g5VHHMZ5pfWNQQp7lSa77
nG77FXqG+YU2qBLv94wyulT7viFcj4oh1CETMV6vuZixmhzle5ylCoAnvh4Hs7BqL5I/paL/+/MF
Oa3MrBehwP5U+LhX/ZA30kGZB284potXsylNKKuIn/KjtjM+iz7RV9kGHsxWTIIdNy8ia8apAW3/
OMlVbniXwmFvmWrvCjseEU7eb0wh4pbg7O8SMtx1PhcIa1ziZbXliakBFXt0SI3L8lRMlRcTQOoa
FFpLuG/CTIAWlinEGTIRuWWaTsvSQfGhaZT56sFTbMd1vlTXpQGMV8Dk4L6wkvG/e1q9zkV8yLAZ
aKsmckRx4o+lCL0xARhdqVdGMs+UaCv80k93EUG2k4+z7jrIEhDBHnJjajSl+1j4AMAqw+O02SrJ
hOiljpB+fjFFMm0VC8jm5Q38nP8uQrrJgfhkVYiI9g8XQUO2Xhpf4bPiXrjEyMFVxjpoRGQ1prZm
B7fhZowiXxaE+GD0tDprgiar91E6vc1rVwyVZMXT918izMIG80/7c7B8A3J3R0XVq1W1YPng7NHM
tiY+GxumBDaXl7F4hVzlnmeMNMYigvF4OZFnGsBW2PnSFkvC1jIwQUX7KFCQmUJ4z07UpgvSOi4m
eEpdQnoPHB3r+4WpYrC5WPQ1z71KXejvZXlolQdeKrbbIqEJhS7UbAi/w+uCv8+oRNnZhx1tmq+u
Kx8U8CbWpVLk8nJ7wPX5qtZDHWKIdrbhfAzHFk8btr++Uu5vZH5hrbrxjiW7D7dMcF6shmdQmRsa
jKANZBr37ndPafQABU+89XL0mdQAU5Yk41S2B0bSWZ+Fvq1AycnqOcKu1tyFGEcCRsS1RyqYqqev
QZjn1BBytiZGhu6yyZeZHBYlL7ENOhHcMKo2y/ks8bbfNihMpPFlNWrqZ+8a9HMh046ZQmRHZbYu
cflNGA8B83xkSL8MUHDLqlqHdDSvB2tVqPDNmhK213ABEUHo2LPWJliO116S2qM/AQxcDcnocnn4
PSgZvYk8rgfLh//S4W7SeklC//NMRFRtgD5rp7ZXMohVOJ6wGcs1KtGRu/hnoEzw5gk/NunNTa1I
vY1xmKfAuDZKHWdAZwnE+/2+7YFDLHiIQhFArnqFCwqHiH/6NiMth55N+W5j/9NW83pLKfxntaOX
Du+hMO80aTz175oYmu40KXqgiBpAa1fDX3UF9LFehgwYPwQheyZ3GVe9seu3FIHiwU3tBRCXed2q
dPGwgmnvcaASdRkdRSGDiF/houruvkfjVG1xBAAamGjzaRzXQV1V6s443imSpiFFw6/vWgR6JKRx
36uwgNgqptMkAMBwPDKN63NhWuLgIxqM2SA0aJMn/neXHAoKmwV57N4uP+Q4vw1+5ikFlOZ45uyf
VK+OThTbjyLAd3uhfoOpBDu2G3w8d6UKSlYq5puyBPdplcv3Aj/BvHDMw0HW2LZi77WZiygEp9wJ
Z9HaUbV23FW2ymbFbnJBahVKua7pIdxSDuPTQx5UTI0edKXFlrs54LXGcXswGxcujJ4xk7IaD1FL
El2/rm2lcfvqDMBic2DowItW1OG507K88aDyMWq3IMxtnu40uqQIMsybvA1AUwv6BArvHOyXBOet
VlV3rt0silSRJOu7osRZhrc9ZGDx3cSFWkWqN/pGWke2pTHs1itYCB1E3EhN2kJrz6z7YXJFDPK+
WIb1hjOofgx9Hej1ilqxjDwYq0CQyPf8n7MuvCtIjwn4Jxfo0X0hrbSLj7vEJzG90dfv3M1oiD2r
ARSFaySyl+jU6VDSzslHeTjhAvy9BAf9aGUz+auttFI9Io75pnueFmn3GNCavX4LsW4q3Iv90VYk
eJosypQk6Ow7ByQpqJ5F7oMvfLRXyQaWRYdbejua7kY6CpLtC59iQCaDzfp0h/yp0lO3vPmGc9wJ
DEOU42xew+EMKTYqx9qLN0aUSf+ARIK+QpKw/b/DUT7EU1K1YL6BBCE6Ss90XJFxLtPPAUxkp6Lc
rVKMsuyo9T2JPF/Pq1k4FbOHvawg0L+TUQXjPaBxGZizlGdWc3+sZ4hYTs39qKubGHE69voCThYB
HHPBDZPqSLpO34dW9X9mvgOOHRbL+sybjBJmUjMboOuyheNEYl8eWJNpjJFsiHNnqdMWvvD2G+va
dBvLjp/f4VmcnRU7WZjQqZbEBivJeHCjz4TFjP4pH1NGG6HlLqvuXhRrIftlzqEp0DzL87ULYFO4
eTYq7SG0ktFzx46xeU7666IdgJkAGHZNkzDcf32VwxVMATFJ+jhrs7n5kgx4l2CWMli4VKie73Ga
DNAJN3G2CXKAshHa/NJWkXRfFkkobp/y//kMgmTMl2BrIqeuC8vKN5GsUCaeYQbsLF5DOOYtyZtY
0gE6FTuS6Hnu03mLN6yNkacqXfg8c3Uq7DDqlZM1F5M0pL25W9kdyDy4+8Ph/eJpPy/poMXVdqD2
+YuJj51AtemTRvHNDGlQTbTZSCrFClhzPWQwdjfNVaejLew+Mq7/vh7K1Mvh28UvjhK46OFnPVxz
5ElulLr9BynsxwQyiY3LZMyV8BvojaL5wWHY/VyEQ0b9b7h8ROReEe0xTFhyGBSkOboZ5IUm1q8i
U8daCvR1j48cSy/ksHhoJkresPU/0sloxR+tlLX9JECTenolSlu2ETa3HfPIQucbDsRYkWZLVTiA
tnS53npDuKQsH6Wii6V3FgoTXUFvlIemPkxnI9VCMkatWvgtiNGBzRWowHsqIv6Hj6fm/J+WQfJ4
Fg1qPE7jTevFs3BIUnAyEquNnXZTl8x6mhGIRNH+3IPZhl8s90VR6A7dwmeG3c8jNw4uZZUuudP4
0HlNOdm5f7RFre/tzzoPG7Rqe2rmeZsdVdDXgkxCcGqZOyz8d8UwwaIbcMusbq4GgVPDRq5sVMKe
tqv8aEWhQ5aIWr6zD3ky1hpWrWa44eOTGigEaj7JY9R88i27aH01mEjgFBOjscbQVkym8W9xERmg
sQ4svsUS0ejJRajAS9pQkgzNRsKYi3+5nAFQiKS4dc5NJNxqhq6K45/IYfgH+upB3i7zUg7T+IAt
RTnMVEkIDeyalZFvWhGgJ9wqORQDfqNcNu8P9uDt2bfve1Kww5IHD3kJPesbOk/L2hpf8L2RQ/U/
abgOHQF43Yb4hhHSPVDubDBo+UNW9M9r5LqnTkBxe56855kPAa2mivIyqpvG/Gv0OCzd8IK0gPWq
bk6eBLZBGzJv5Ck1FOOk4sXqJTUooiIuG7SuAdzl7Z/ioyGnny6OjCEeTK3QUxzqkQdvdhxR9RTo
r8Ku3f7LJluUf+0Z6oB30q567vO5al7/FwjsVsOmKkzJsTLtij7omYHdFNrMjiotNFFIHDdAMq0E
YrpgT9CCWWZ59uDDfN8yT5U4uE5Ns9pyRzvejkEfrahCawXkgdhECQAETy5Kxzu2WQDv3XA9dwxN
bw5b081XCUfbqnL6HcyWTq1fs/zapNCo9uGnZ+itPNGWSB+NApyyaDkup2NbcIr79RN/s7VwA4rG
yyTbyfB0DAswrEjvOST8nXNoRzy//TW5hj/tt1CsTi9KyiSK2DXYE3XpMkIB3/X6hzoTMLkG332x
ohoUKonoNB5nbBaoYo9mb/gF4UbAdyiVof0iTI6RPuW84z6mDSD0rf5uJH8lPAV715CHHTnzFIv1
RzwSyZRaXA2JEc4TQYdg1p7xag2caF+YeOUqso9QMAFp9Fl1/qd4BJnoRlwfjhi1AEx9QjrQNHn2
T2GGXeNJnytRDVD99xfVxcfEe/5mEWPaNbPiJ0uZsne+qIJ8lKCWxnFaaPW25tiOZZKfoaR4B60v
wS9KUuU2OTREJPV78rdnENAau9ksGkCwWfWs/7IocursCIOmiJ1txjHyfHxudj4LlgYoiT9ULNPn
3lRIxEuXeklVlzJvy4+1AwgRaM9RsJJQhejEhM1LpwNIPnsziBGP8u7Kezc9QRT1z8SR7DAb5fpQ
hhyxlNLXOSBSv/qEbVHL4clj8pLQtODIq6T5WvgQO0KnZ0LxE/XeQduVabMkaUjXOm9JGu09bCtS
jUDMvC1vmtzHz+YrhE+6RlPE/oJC6k2GW6ZgLuo+PvFwecxRJaHGxv0zpKPlq1Ffdr/xIezmqekL
pdRCPEUhb3VHIXGCq2K52ca7KTgk/da6PmsbpV+Z6kb1lAvAGdD7U4JjpWrmgk/NTgdL5XlMHSSG
5wVYobQup4fWLq54x0BX1ORqVRrjXv51lwNbYXfHSbEHqptl3VcEiGV3MjFHNqRqrkVH9cfL48JB
v4S+IOZp3HLJr1yXSLBLSEBrvDTEzSBFCJyfFKwKZF7VgDOiOdUd5WesVXTYJWOZjThcu8N8vhah
TNuBM5kbyEdPi4wdRhLvz/bN2+eSJtuEImRo8l16+ci3yb17uNeHQvyKdhpp3GdCa5MCgAOISIja
4kR9arM5Jolsoze6SWwNsAGY8IKOS44CEyIxVmRSKFTzPJihND+ALvq/C9A2EjYnY3dIFSw5yPJp
MCCicQQJvCClKvUOAjzZYyT7cM08wmd4A+IlUcXxzYZ1ZWBu/n4778tP69SpUcW7c24FRVgQfrwP
joIEvN/9bPp+mSczpTvCJRJFB9/xbJmil80AFZlMDiOyEAEgqNhWoM6cpC6u9nAOPOXorvTIYxbh
0FCdbe/ZH/NA8zNR18JhFwV30hPzJQ7LVgiBVK5pem3aI8947YivPVmiN38MC59tOUqMpvdQuN6d
usFNcsP32YMhduXs/TMPEEBv3pknMrl/35rOCMgEHPF9KJs8A1Skmk3sRq8S9G5TKhroz3uoihhq
zjT5YbG2AFDA1bVeNj4UG2z8ox5qDE/LEi2DVJvqJIMWqnxD85s6qYSuJgNl9M2q0Ai3rQYub6uP
AYb2Zj1RI8AsYTO9PhQzrzFiUW+n2Hm8Zj9eO34gYXxQL5400X4aWiGn6dzV5VYQn0zeo16/MNxi
vdnFOEbn0Z2GURUgAUMYbHSrzE8+fAAFlLeNthwTXAJL+4PsFi7ui2uiNTw4h3dXksdHnYmBGIN5
kqTzA8L0TZg4RRA7wlE9POdl30kQ/TsU3n8E1JOLrFaUO8a3n86stXJwO7PQQXSceeIhC1keZZVX
LtQuVseMQh+ZMPZuGVR+Z9kXpQ8OOzS6mmTuJy87HW0XKx+LU0NFpV+l8R9PI5jMvo/2cUrACwNO
j8kcM1Ud+SGpWlYi3PAGliHzN75yYEP9YCs3SAzcO/t28o/85C6iNBL/WAt00TbdnlyjTez+3yXz
JyaRCrjHMejArD6cQ6cGCTzTQRgfkWEXkqXxFADm4TweuQ20+zH14+p22qGH8ZKW9VNsVkNUHlE+
DGz6k+80AsVdalzV8tzWA1au6A2sUSz+vQmaV7XHtab7qCdTdF0dCFaDIFEEkfdYERBjoMrZR79d
OravRwdDJjSTTQpTvYaJz7UJ1H29J1LIv7tJUqSaWeDInQKPT3f6WjVDBNH+D4D1vScWRdCvUH6y
GbtYQwCy5+rtTHdp5uym6EDIMqASvr65b82z7xkKyRtcKCx2bw7wSBBUrx2lW9RWTvIOKvJmBFlG
bQKgVSbZidQnXn+z+0GzCc/LM0XjxeNMSodzDa+lKZPtIOaJZcif5P1akDLK3snbVgADPvFE3G8U
I2uXfLDbU93bxT7IoTge0j8EfJyZoeyyqroY+FgR2193AwUxjefpyYte17o6Gox4Ip1awvGudQ8S
4UlQjK/ENroXho+WdN7q5JXVZuw+yFhjbM466nNpwq+CHcRdKNT+i693i5kIJdHu5DqNpksAnLEg
L3WZ655bOq+pwkNq/PplZK2httBrSphun09DphzJ7n2a4OkWq68AVggy/SNbxx0NRxhzezFqEf4e
oYnetPXKCHeuBgUKhglrlBTsDK0CnN0dThCilGYf8W58PllBJwQ7kBj2F4NKXsX3deolXkewgSBZ
yFmBDQvqAnHGUlX8rtTy6OFPQTvy1QciKEnI84aphjrJnmnDK3Ylb3pLgOO+oUc/QHlXQHXu+zMA
JW+29MdrZUMMtjbOFu/ZElnzf3qYs36ZXedTq1gqx8AT+UzgbNPDaopsmkFy1moP8bi39MnrNd/8
fyVVE2BzjeteII4iWAxio1L1xrdBm23H88ThalfUC/q4p1ALYerbPMoTJvJHziYzv9RA3hmo4DWY
WsMUFnYNRD+J/qP3Q/FgqMsJnPnMhYfaVATppyyui1nyhbp9b2CvbZdZz4kioI/NvqReV74dhYHf
bSOeMv+VtIzqMrm/260iOJVzt/1AqKfHbeLVY5AnOlG7kkAP6L1hCiup0cLNiwr1oow9tQ9TODE/
K9+aJ/ZQuBbxRK6uLw9RlqzUykz3e5Wm9suYX2s2mEJ/CmXP3SVZZMwEhs8u/+Skn1D/vac6LcY3
kbReveamXEQD4eYGBZR1MXvHs6Y7M3UUEIbxA/0PCfeJyzx9U5kV3sL+2OqQGX0xQ2oEmZD8Mc6w
IUYDu0hItdCOq4c/Bsiy1zhXAPxJGAGFAg3BK1E20oNUJi5OZgOEKvhcW0pHBrYIiQVSnDFU8lJ5
dmq6Y/2hY3BG0j36d4JEvJwtC0OVE7bdDvEGLRDLFf65JNuYUqK+rSJKq6ipRZL27LruyIvwL+fH
0ORTT1O7gSY/RH3LZZK5K9/siQWIA+BgHFJD3lir83+vhIQV2UrLqaue8N6Wea4XjkvDltwrt1dr
SNbru1MpdAcZYzoOcM0wkOzgQOSAgYNfzCUVnCXfLPBfhXfxjaaYX6/AvlNzuaa4nLZmKUuNQNj3
nlQPX8o8VsKmK9wRzcf+7g1nglcYnB1JMcwoTzFEZI4yMtT5ExoPsMSjGOxTR+65jhl2sbi/iZy4
CbKqYZxDZb1EWO/JGHdPmEgZHJw3V7v67HCdk8Ee3LxPVGdQFFriUCuWJIPanIvqP0Mvq87Lm5uw
VDJvEbi5D/oNBIHLUx3E7/MEwf+/M1Dfjf27Di7I2GFYazLtuFjuA5xuRQi0znpg7SDMtzlRbCZL
6/qxVArqQI7aF1GE+CHQSjw3YZNfFJQs0nAbu+e1MC+E+GkJERjH8S8JDamTc0ZbuVrARBZGga5G
HaRgfJbqdDmjlKrr5vegbzSoNyeFyqSfvty5vPWQa+k1mkPe65sK5+aeUh3dLamc7n/8lNhfHcnk
Tyli5YRBdjR/Q4QXo6jE+LoKeX85qVmBPzL7bWTNQteHe6ExyYw8T+ajgkNz68/fzqfWZFU+ppO+
PQUKXEo6IHMpZudi2dDnkpe7HGeFGpQckHE8O/0hLvCztmErLoQ4wKDl2CAPnzcQ7vPDFQcAHupk
Qm/NtuPURoP2ngvED28DbBjotLA77B9gk21Zve1C6JdacHzkRA40drowp6Kgzzg0i6fTexZ4XOaU
XezjnJaz5Ve84r0la8dvHM3mNCK0LUg8QjBU1xwcuIDZ/0UoiHlM/FAlEoqIlphPloAC4n5NsLaR
S02RIg+zXtsoEgUyapzKd6ybMnYml3aHe6M+SkERMo5vP3sobMcBrZmdtHL0iE688+JC5VEFUQFY
SxbYON679ou9T9KOJebmUbG5+4Et4iUlBHOSQ9BxxMfI0582nSJ6WMpubl76uN7tr9wbqBDe/4JN
WzQLORbk3Cuq195AiHmDYXwdbV2v5zqne6FQ6NzqGKhTAWsdTL4fug2Crb6QwU/ffkFbNa9jO+Jt
mumh0Jp3PhZIMa9IDFz05kQGSab22wrDxYUfHlOjS/GDNODyqXVV4ggTJwMrWY8SuSVqpu2bo84r
eZqtt4YwnBS2nxuMMz5EtKdhSAz400yd5qcUQWCvbd56SoyYl4lId+kyodRd1Pm5pRCdB/OWLrBi
BVNzBGyaBmkDDplIBLLbp6z7m2HtcZuq+gJSHQnLRUVu3G9VJhzs4rqFOUXaOicOD7HhyXgLaL1Y
EcUAB8teZ4vZCa7o8zUOmkcK6ymIFvVxKs+NuoTWU/dxfZvNlX610h7X9FXWkw13EIJfQtGODuag
bOIzdhmwbXYgkD5fkztL3C9X++c1D8SAzaoIEFDCr6gWEo+IxJQ28UKlwlr81vep/+1F1+aWt5Fd
KEIfyIPpFA3Rm8OtDup1oihvWrmA0Eo5xVN/WWBTfSTjSp3t3YvljnyaUmLLe7kA/09IeRVshvSB
ZT6r1HL20t3l0PB+9rhKGXb+lgxO33eEDXI7hIN4pg4AZz8Ty7PdKVsFfBq1+6TiOrsz8OVMCze0
/q1S5plm+YOR6xGE6zaHWN4YeCbKx42ODbD3298EuxwnOED2YnHDAQ+KLg3/8M5SeyY6R5MKX1IM
rLjmgV3g6xf/d36q02srwThar+RGJcoVGHHCb8c1Sg0d0I+LwvzIg9NGncsNLXMdJey4H1hg7ttI
BSQtcr/Jt2II9J/3RRtXePWN6iN2YLISxJOUY+UOhKZGI3gB9GNsvslekSetNPWv3pljORFPaarV
/wchm/OXU0s1Rvrf0QyBNBmeA0SRDobIb2uGlLwg4xsAuBlmNwCv2SIg1kbpjYj3HtG/otOnOVHL
Z5rJKmHSlrLSi8NgX5EkwO6zmTml8M/+SxR02Av3kbaA5+4bt2ZgtfSfohe5OQs8D4zBnFdODw88
GdqnjmLbIg+I8BiH2n+vZxmU7tFpg80S0H9VVplmTNm/86anNN5QsEvo1G+H9NXIZHO9YbkfM2R+
iMqHoCnobAZUxedx/O3qFK+Rzppiy+t8mjbjeojzyK+fxjsZUidtIaCrji6IHfAsNKptrysLGr7f
U+a2mF2YhGgOdmxQTZ9MqnHSH35vFbX3jn23sWqkmji8sBlFgWEFxCq/zAPsXu+LT43WNHXTdh+2
omsewCNLvUSX2hgr3iJetlDg1YijyWOVTgS5PIEYLhgN9mbeKFKyfBEY+bJAlgoEcy3B74M/oG2j
wDXBY+LFn9DYxCQbbTdBo2Tiwrp6Oh754YON8YvmLNLyqMfKGKZvVRsrY9xrdK+BhQIbzT7Yxz8Z
wmOJNEVG9rJ4r9FJk+hBZBI/Z5XhytTPA71SfDtQ3pQYnSo9hQ11gT/Cr5uxw/bk9sZvGIVBtuLc
6WIjzeAMXbBu/qCUkKOa08W0eKxPMublnIyFqjXBmAf9mcQb0gfaFDI+AjcY49Nmac3zDyGZZpch
mMDllQG0iM01DYFEdeo9Rmj1BkDje0cObisW2riNPSbwmvgLikW3xe4AUYWzPU5KjFFg1DdTEmbc
mdItRCv0EBNVWnpI47m4cD2eyoAAGbXjGmFyQyt3OEaXCS+aycM/8mfsIoijFT2foJBoSRrV4G74
a5EGfJQZ4eLGZOT69eipn6yQCqTWtdyBmN13K2Byv644wbliWtc2ErGNmsmoUgeSjCekTPtJkq6q
cCKZ2hhCF3Pd4IkCsM8ZTRIT9KJmaSa51PGPFn66duH6TRMYn5qY0/AV+a6+GT7erQXtq1JrvwM8
OwM18/bAraCSf7nPN1dDc6guqIV8e1deUgJxCsJQDkTTV5jSYIcLLfc72KR0+gcrxPgDUH9ZIXr1
1NqKBhMiZSYmG+B9n+GcpJA2RCzM1IDIHtqLhC+JaoGNkkRmoqOe00e+o8cs9RivgdA0bvyWi8CB
qOkxryTCq0EIl68kTCQFuNKt+4ErOP5LOxqYpqm6Zj7wFisvXa8eK14u+bc6l9cnVxCPaV84169u
JgguUOQ9X1zgo+vww9PdPVAB7cmqU1eVZypW/wc3f5+i+/feF9u0yPDkBS9YJH60+LGKD82kEfti
T9DM0ZwkZBfvsnp3IecKlISe6pyYyXrqv+XP3IA1nafTKb2rYVpgUexU6DFUyXI2CrYNf0Su3ahy
L3Sv9RG77zwlwDeWiMFQ2so2Z+ODUX+2GsF3JkkozNJv0RL9ebFV5BHOUGkzg3p1nm0BzWr8diUs
Na93O+yvRoXgAaybY+CIPc6LoScHMaNT6f4MVqvuN8ipRSCWyo40+ptWJK5iMiQri4s4ARrQvo5B
PXHcjN9r7LKJW2hpd9vcrYwr8hxrZdEEWYxHh08wf8hIUonpfdmgGFUg0rFeSzS6KFuPeKXRSnvO
zXxVhsOmdl1EzLejcgrz8r6g/Y52UJ1H2iHEz48nWj7YFNMiDA8FbroZ7uWfEp3fE7nqEr5vQ+QR
oxSgiuBjg2VGv4jmtK7oCiTjurU2wDR/uPxbBG67SsrFmIx1xucSC6ZyiQmYm8465JQkTqLGMwk6
VhgLmiWAsFUYSvCEvI1HeJq1CYKsKwYWP8GSMd1tFU9kAys5UeUrBh0ct3RTK4uag9q8AVxr9MBF
DJA++Z3Uk81hEz9Zt/D+WjBkNmAnVc7fXw0PDMiOgY0z6J5kDpPv8el6ucapA2X9Dt3SHy+j6F6W
wICJ0iadfrUdMbPUTiGU1ImpsbbFwTCZqn3LsWq4uzQly9FZEVcjOz83P6lfZ4LhAXIq/A9b11A2
t4lmZJ3YeOjsELLHt/XG7TOQj43ShnoDdRxXfFCbiwxW0GjUNnhVGeaYeeM67DzIYlQKVf+jUds0
5AEObWPkRggNF+Tz+fQc/CJ2fHLmo5CGH3jSvp1tEGXst/+UMUDUNXyv8qEgQu5Y/+56p7poqeUi
x6ffslF3O3JJ4ze1BHIhJQfdz6Cr2obzMLntvSrN1Wekezhh/0ZhwUEIbwgfW7z5//hJ0HaL9txS
SpPu0VxWOB/3qgkeI7fnUmmpVpg5ZiYqwI0m6bMHiTfQq2ZAgdlGyQcJB/O897CvPcrKtkXp1F+3
yOEMBtfGS13Q9qQqPboWnor3dHxgOzdYk9oEluDvscAYsYEFhMN7ATp8QdbWwtEwJ+d465DF8gDu
jabzjnUFGfu5gF63EKusgGfhQ6SD/0AYo9VbAgbjOXgkvTS3dY1LTf8FLvJsYSC+pYYXGRl/39R+
nlFKfo1eGoQGKealBuapzIU2XdwmbB39Y2E5zZMXdvJQCUaJE9QmXJH92O7YuZBTU0qEOU3sUkWi
HCaQsHA2lzwmwyjeXxwUFe+A5P7P4g3SixFpfdeIr06PpyJzYMAtlqvNW6EMnEeJFNfMQxJKFNSJ
WCEKGu27bsk3PNAwu8qpbHOzRYLXTGbK+Lgq6gn+KTUz6UtS27o5GbsqZKLvjpHvCAHyXV6JtSZ+
eJFDcBaK/1m5gBCdQ13o3oZy+eIzbJ9tLDEhZMKeX8zZA0ZNEQr0Bt5QTf8M80ryGhfT6H5kGOlz
K/mUytpbHSsnf2mORM8Wz+NGKDlJHqWpypjQjcQl52EBH72NcV30dy1w+GPlniQJ4qjMd3mhs0UN
YfP83tILx9YLa7YlvLB3xYRr2qSAPoRERBseh3J9pNdpebpi73g68+2u8viSZe6952JvZbWQZ11d
PYrHu/LhslJ+Q8Kx84wfNfWiHQv6kaJP+3C48jf3qdvSLMYSNqbvFTOe5nTr6lUKfdi3c6qHTwKY
b9WXmTg02deoKpuC1LtaNWiEtserspunXgqpbVN5AG01/j17IpAndfQGMxpDCKFUDi3/OHecPHVr
bXKViLTqklCpuA6h8tDVkhxwCqOVjq5QNZd8CG97nUl/3r4DXoIS+IS3heZaCJ0ejFyXii7U9KnT
r1wuGavpCpHvmAtbriDPQY4GfGu80U8xBTnXJT4iiPzL+fT1ofQX/7g8YxpUjITcQABFQMBk3GPz
k0RplVa7+GQYbNh6YPOvneNIMaqKYv7X7CqEXOmMUHdHK77R7QpE3KQWKiJqglGDsjV3XLPs2Clu
d2jfdXADppjRgQGj9tIt2Ao30R+5htKRB9n5wHD40euft6IWAfA5xaud6ls4dQaOrhfa753CkDwO
v33/5wKm0jI9pAMn9de5Fkyve8M5Id52609KHTVZNMjYbcA3SBy6mD5SXzVWwAOET7ozgWU8aAqy
7bnNVkX9uw+gnj7J0Lh5Wr1NNenv+WKVh8COH1SgYJ6VKIiwwBECNv48IiLC62xWJ0kwR5Wc3Vx/
ADYMCidm4XsxudJQWjv/i7hjGKeoCo8TY3P/mJ4yFF63RmQHKtapydolRezBD5S1aw7VYFg3qiXQ
0Hk5b2Ggxpo+CVpDWJ28MXN/2CZQoEcfVrOod3ckF3TX9XsFuudUtakDt8bkpEi69Gd8HR2sAbl3
tNYiqvE9lNFIXw4oODyPhWM4GTU4fCkVgNhuNiomNX5s8k1meDNaF54rV9mpEPFU2t0SN07fQFlR
eHgwyWiOVJ10+tVNKdrASyEHD+ROQcbDZ75+NI6B+EQ2DeTpPYxi+TyWmcvallVkysO4G0cbFGOL
mlb6qoXvb8cDDalFX+kTzkkkHGzDlM+UbvD9+/thVJvMZAogJdnmJ+6947xX/rLHDDuQktWMQJyE
0x4yySHH+CTR8k5Lx6tNbCx85181CNWvepDOiyBBM3bs6AnWUmAIdNYfAFaZukGTTOjuuACNIWjJ
lgNpIZ4X9b2O2RtmZBiuzAbRCZVNfJUqMJ2jZcvm5QoMNfvuT599n1yx42fp07vdtPe5HDIaSEW8
G/YqX0eERnjXRwo50KM/6HX8V+pmxZCx2qTNH1RlMwhVTL98t9y0IIn3uUuophmIgAIfOPibI923
KEsYd4vM8DgA/UhnSd6ZixAwZaRmtVW2E6ydF4oUkKGSRInRFm3npmrj4RSyWWd44X0p/bTm8BGM
3Wh4kypAzeqsUWskHUoDZKuRTfi+goAEtUjWjF/rtt4h7vPY04FuGAmPrHol7SgqKhjH77yXKHHM
UnjIUEkvJ3HmDy0qzXgD8wK/LWEIPEjiYaGAQY9oHQxGwN76b9ecJNiA37RP5Q3xY/DLkPUs+cYY
9oyw2eSRSvBMclyN6yKUKkypL9SQHesXXITyqeNwARoVt7vX6o7SP/967x/UWi/fpOuzcWXKscCU
qrqFtWLMXBngIuVc1snullDmwJIG+AsXMGTF/UY2iQFaP5/x84IaYnA6WSoFm3/tOLfxrF4B4Cmd
nS8mlT4b6PBKXzq/q+q5/cufftj9kzB7hDe8WqOXDOHwWBOrmnAjsSJDjyeqMGAbk/UXiuq7gqI/
ZTA6jqnCAJbO5oDuilCAYh0wBjzyzX45c+aK+eGz0216VwK2U9jCUQznJ4Ie1gpNdruZ6oPEnHfn
Wkihs62JV++kTwUnllxAoKUBKQxny4opU4MboM62FI+x54vJAey1OIq89mcH0Jnr3upjZyTxyfqK
0mFP1lXD2jhg+DqcswIc4m5au1/SCOcUbdrfAbAkxXGIFucxi5oj3jKgeiyddGRpTax7PPAPn7xI
V+20T84KlfdcDu4mkusTlKDv3D10fOkO8f6aQOmH1hRfiuCFVRoS0YYXXTDhxfGDYB/Ekj5d6r/M
rgmmeFGxD7oGV6fWuyAPMrn27LC3urofkmB16UZ9yz53bA9neQfnEY44bYtxFccXjUpQvzPkz8kM
jecffhBFBjmcPaz2tSev6RtNRzOSTnGqKLDdDuAt5Cz87hWqyj57Jr+8A7bDAzbNAIQ91+2MCXYe
TeMMhUeTwOfkzX3ZBBX8vTF/V/dx/Qo3JYG2+zJBl5nISaC2IbJ4m3Yo35h471Z+nG+6sYQzU7tn
hECUoS0SeTPQ2a0SZCTBPg02U3x6ymWHUEtMuVcKnWgJ6KcRYl12Hq9crOxGBudm2g3lJDYaf0Ep
h/PhqSOTsRhNNnBybizrWtd7dJXCbpFFBcWGVHzpJO9EsTFPbzqWYHKkePSt7HwW+fQxO3l9XvPa
tiYt6STe+ED5e/1OMeQ8DG4Xq5xwoyLuGB8Enlns2E7Lgqw+Z+qvHkfvKTkOFPtfwCTnXIgEa2zh
jIl6HJXWJwmMozXQKYxfZhPT8ZyIWoccOxc9I759/9aJbUAkvd0R8gAahB6fTrMCslkyR291sPuS
V9Itf0+5e+efHGzjQizEWbAPXKrB0dyi37Ti0GfcwsA04e5aDq1e2Hg0zTSfXQAwqE+4w9G5Y/Bb
W9RhLTxINJCgaSdNYy1C5Q1ZS8JAP/7FvmMNB1QdChJEOJcD3HBfnVhGUbONId0rvkEJFjLJjpdV
DOQc7sIfvioNEpc4oVgSlJEU1A4VMOTcZi4CIocwgROUG064gmWbGxYo1lSUuzOZP666qij6up9h
bZleAiObdFT/iELpAb21GkUeoJJqj0a6wvIY1W+xaoB9UmlcVLPUM5Fn8JtxPaLUAPfG0a6bj3rl
bCLYeDUfhtXPhwjvaTaewaEO1jsuYJrPLXfgcx3VOnkEsLoYo+Uk/bQLPAexpRRrnFavfd8h7NfW
+IoNJVXiFkVMoZXNoDzWATWNvS/fDZ5UjZILhg2Hbj87BV40WJYuaw0SeFrpGF8X0cAgQoYzRI2D
KYWYph/8QTgKIhS08JJ7lwqXBXgpe+1W/Cut2Y2YbOuasQGr6B1JSNppcLCkqpkOh3gg/TXgB72c
b8aRT4xxTC1Yd1++I4wiwGLghJvf97MkEBlkePI/y4GcTHDadsHx0GBGtf2v/v8bIoc9gUEwptlq
ygvv1iExGGr/SwE7I7Sgb/Gi/tEVNOd79S3KHNlety57aPki9woHIFyU0mOELgR+bmaKRCH0NoOj
vitB0gD12pWfhCjI4fsvX4E67gmumEm1qWdyq7r4yC12pxriPMrxIoBBGHyLQIRXiYS2bkVz6s6p
BnHyCXydbhOSBdbJjDd8f6kbQAn+sGNXnMaewnf+QjwRTWRSZHELCwUjIqe3cxh53FsiTnFlPoEI
UXhb/CDt05WPAfJcI/8kI1o4hzxoCEDmyPKaliRKtIX+FG1I+FYOlSPWQZSq2xhhn5OOldUDvxcZ
OxRZRP6dbltI3atsPuTLUQPePCozoxXOHUZC+s4fhok1ZCXE/18uEdG38NLcjahwpZcFN/K7bte9
eFY2XivF5nl0/n+BI6SftRxzLFReFNts04RN8PhtvkIW1R71sdbTDB++8IhDI7pkIMouCV374vWx
4HlrXhKwBqalD6EltkMo0xXitZNrpJ0cs+kJuTOLgyg0ySieF0Lp3SYZrbBotCVsaoovTt+l8Y7e
/JjnRdfzMtrrOZV3XGfTvmy8TWNZoLxL4RGr+XhyTPG3V8wXtaja8V3eveXcKZ8762GkizsRweI3
xuc7kDyhkFv5gk3RYzrGwvzDkADJY4Bt7SDc6ZmGZQOtwrT4fMuuRjkIZvon3DGKczKIRCh5NmLy
OZivmcDlkEGqqpqiVolwuayqZrQKRVM8Yqsv+KRIa9mGwn/xkA7koqxD95ppIvZJN2gvvFCnxJA2
K5DWp39xA+AQlG/edNMrkz3V+QARsi/fiE0cc45kVyXrugO9oICQ3IQoTlW3ybRiIjzmaQ+5o8xV
6kI0U+Etn8w1hh72d4MOwhyRj8aSqbXCM5/TP+VnCMbTat94B777s8twol8FyRA5+4EWpsZmBOOi
C5IeAnqc0ZOpaA72Uted8NLxHBBrZHVoanMNZP4htPC7fQ3S7DyyhsZkua/mEMEuV7Z3x/gFipx+
0Fk8rlwwc4PrbGBpbuXqKJs/NArZmSA5gLp5DMfxX/09iQVm9g6q/YltCpEEQjcmoC1Dc6KykkHT
kRaST/tXIX0Hi3fdAWbAx5O848QPIC0+lrEkaIpNjNGQuwTicUJFuTX3i/C4k3RzM8Oqaynf15wu
dav98lv0iv56FxqUVn6QcqaRKBcY2qEq++qqBTEGvR08RHmHYBtyjxuUUqtT2KDbXYmcwZcG+wQT
px+mdQI3lVt+TswArea7MMpXbRnK6GI7Trfi0evPTyvUpv9bRobrNToV9MVYM1nIUX5qktSwkYt0
K3sMf7wfrpaMQrgActPLJ0q566fL8L0mSCd7Swn3EZvS6xTfPPgCH0Ah5M5r1+HWFa6LK35n4+B0
4bsYYCLrL49xRkZjHlGWGMlQ6nlZ1zQv2aPV4lRLF5Jt/sU07emwv2+ruDFedyWth6xqo07EFUm6
1npVF+UWv9TvCzwU1TGjV0skcsydt6nl+/AChJoTGgReeg/ynIF6cmIp8RVS7pmWK9j9m4ZR3l2i
6+Kjrbp95ezdkBTus/78rzto76mtNtvlqEA+4+yuoLeSeb0fnb+2wiDb3tfkibm1CSs4FEc/aod1
ggke4R95/5YrLymGsHvXhDIevK8jJVVCwx8iu6fCtgSoG0cRPsdISg2Mkif3ZNYthMKPs+d93woQ
cE+cY7ktq4nlAU9W2RuuNEIwUbZy3BQ1m3br+ay1TZfvnU3PsW3qipJMJFZw+jjhQSTI5pALDdOQ
lckTX2kr9LGqKeubpxZTP6m95IxjO09EdhgCK1BmZ+ClmiIyl0K73PFEIa5fAjsEJqdljWaBlEgS
GlFGv/26/65npXZ/e9EYqLlFXdg6bms/JwNHCViRZ3M+5e+Hxz/Vag2N9Xc3vGjLlaMG8gYaoQ5s
aqBkiLKvzeL5uX3L4QXb1nfUCQgdKFqC4D+VYagk6rzW1gGMANvC1z0c3hg1lEH7J7zT3YKFfeVW
06Uq4MdsNJllu/b4z/o9x05J771Nd6YYJSPpwngvxBg1z4zXY5xxBnGZM3HuVMUKpwovaNfQj+He
s6W2qLzNzhPBKIPabhgbCGLwdxudWGN4YTCMzEV96IxdHW2bF/gYjseE+po80nsb1ITMf5eyZDgh
snpm4Nv4eiBK5cGqQqCRul7xdzz6BrDCfwRlmB0EZhYXZPOWW4IEqH8x6jueRujuCF73IGBZkFUt
VaIuGclpwO7o/HxkK+PZ9OH7v/RtaTfgRdmOaOpQtl+7duaPWJwynnDx9mPZiHe3W0GjPLw7MmjY
yEupobLLh7HbxK8Sxz74mpiGZG2ve82PhGIVtknzfbIun7FRar64Tvevql8667+4SafX33Tn0xy3
y+QumRyKzQhZuXo6xEDc6BivKKqJ2DjM9Hx0b5C94csQv2ozWiR8Ht+LHRenAGvZrQ47HP5T+vdN
trKzm03z0WYQQS6EZ4vw6OoquZ2edDQbTD8tRBvxenTlCQGvD2/3T/zPkQidgEEiEc0Gbb9WCat3
6lN4EmGv2zKtIhTeFRAKdC7fY+/PHfjMseFPJaW+kZcSlJD4CnILMV5hsSHQZGN/wMZjod8jHhsi
RclZSbT9kJGx6aY3H+pHMo+bjuEeFHTHZTOCAFkPJs2BqUWNUNV4+G5C7yy1ogDulXLw/t7dj7eZ
2sPrzl9WRHGnA12M+fMXsoxA46jh3mDchi+C0thuMsnK9gVWj065Ye+EV5VIE1bLnrU87ia4V8cc
voEsI6WpaDK6BTf4l4KYj3TZzMIMfrSP3TxyH2OblRXK91A2GzwXkll55HOamOemBl/Nvh/51J/0
dKDZNmt1jxVFhMlaE7GWPtjl6zUrqdilMOy2ctzTvC8Pv79WR8UJuNwQjQRl2E4S/pjMZZkuvVM0
JwuDXgdiEXlayaIUxmf42mcQUz3RGNIF1XkRPc1UNvr+IUUo7LIvvLZVXhaMN96MK4m9VPpAtFeM
gs/LPWB/h86beJozmWX7djPcF5xzRbjLIvAzPAj5epAioY/p8U4lxj075367p7QFXh8htWVLiSz7
5f+ooYJxwZ95VYQakXQvO6bhlgL9kYbskTsIRGnDjJay3wmG0GmziVcrR2/zL1mDiUQHzdSamFv6
39PBuV/0r0S+z2P8bC0zPoCOWt9l+typzRrh+ID3DvvgiPtAoyb9hH6p1Mz50sWsG+0I5U/1r40D
rCs3A9f28lbRd4QXiCvPvfwzMEWzI6whNnE/m+gS3LLbfxbpD0wrWZ22Ci1ccoK+BPp4aAyWoeId
7plRArRCaGKor3Y+p0cFONDnbg3y5k8rKP3rT1u1deKa+QTwC0VYjFbhXEU+iJChTx1ohPUfq3rJ
jcPTrFM4fOlDwvl46c9Rzlcmg6Y+oTz+oT84RaY/5okldvg2NtXxKSrW5bcYSTPpHJpOliUH8O6r
0AaN+PduP74M/6XsFBGRO+fRt032BqDIhZCPribLqgxs2Cjq0QuHv5WlgxBccnu7NL/uYQ63gv+L
pzLPcBNM5Ir6BPa9ZIE96p+wuWHaa790Wn/Oh8SxpjKERMpZP1ktY7D/JPXzMEfaTP8Kj0m6HVm7
D1Gte1lB2VKTfL+5wDSxjIkE+HAfLOUqPzmEgBFZmqo1H+IbrskYRp66bAZagOhZ37x1gctDV8Kx
TPOgqOHuOQ4LtP1Y8iM7EFpM5bdQL/O7hqSOLrd8G6oUXldY0Cn8FYud4UM4O/Kb3p8KXXmvQ4fa
XSNbNy3KokxkZ/V2kcAoHFZ9ZzJmTbSacejsSeVtqCa7oQsm8P4m1+BcoZ63ML8Day0We5/pO1C8
WCGiDxFSwRUWfmtdqbBiO/Afc/93M8Pa3KS/e+pwfPMI80PVVLjgCg7Yd2kz31VtvQy+dZdvtWD0
NtsO4B+dt2BI0O+q6+OiRZnB4imBK3x/WSVQHtEb/xOHuvpvIKjGrpWy9MGIqdDQtKHVSwTZuMYV
b6wVfsrWmazXNqHggSUBRHvQQ95NuUaf9udnVr14B04RMOLKhP4lqqLwGQcxsiUIWpNKZfsIoIeq
nMeK8AVnVkJc72mnu2Oa46jvW1iLBZ4yAzXDwGzcWfqKvmp4vqkFtl0pPO7jX1h+txFl1TMJ9egK
ZbF28OOf9IV0+LAk2vmO5suZ5cBSm00h2v7O7cHw6pBlmKjEON2xYSn2AgVnNOelLdkWS5riuxF7
z7Zp6P0E4Aeh7mlKZm27oo5AZx/riusiW/ucn7EpNrKnrZWCT5UIfKd5oAH/DiRV1p5waCBJXsFi
OitvTTkkzgZEWqTXbGQz0rm2ZfGijsAIu38V/42YN0kVEgJWoiFgFmK60P0miQAudnKQNZkMc3oX
e/TSMy3KQ8PblAhiNLhCy8cLbNCIaIlUfeLDI6ax14f02kxLJ8qeHMXUuaofbgYRgIHBphHEOiCz
qIJbLjk6vmta/+mp8upZsLVNvpViPCBgeuWby82s48wOJZ7YcLugKM5Jx8KueGkHZE2Ds4O1Bqqo
MFMvf5tQM3Mlha8Cch8hxJYqUYvV21EuAWL6DutSZ0hgR+dgqQkLSAHIOYDg7zugbmB46PlHqD1r
PCU0FDO8bUpq2o2mXZQ5wp8DF0m5Ojzr740mUnRTMh/BMSzmEiJ60oIOXoqeKi8E4ZqnMofaRqf5
IERGDtFMPXCgLusQDHQt7kFsWKNF0wg38w2MW1Wcp022pI0znEHLE3jPF/QwvJmA+P6qAHI5dXii
XEzS77Y6SawtwBnmO3dcIFrDvlpACPikGyDh4GN/hajAxaMlrk897rIViSIdUxGwhCheIl10xVz8
Brn+jke66qJS1AtKxSZudnzfqyD/CU8HmyU7VpHKCV3vQs1hw7xTZYOPwd/DCyXtENH90NEJ5+Ic
uV7AP+wgvx/9iwqILJ6sRUMdSwiUDSNtBcaTCeglW6pGSEtp+r6K18fDhTuHmyVE97+yCP7l7JO4
Gas5yIPEWrr3aZEW3+NfqTDxKbKJur8eTnUNFWYrxLYZniQXjWvOH/jj3tgaJ5x5YVP6QEbSmAnN
Tt872trehm0ToOL3/Gv1uldmF5EYWJY9AkhM1HHcWSLoEk7aDPuTDi8+mkVf8M0/MRfP3mZ3zRcO
YL+jfbHW7nSbRM29IZ9GjN1GXvnlc2uStbvUi1sVxGHtgk0bcbbFBJ2BP8KOkRx1R4D0HDXcWOgV
zzPs4qTrtaGiCZU1CSS8A45N90llTrhS/xBNPhbCP1yJ7AKLiHJSBfNhOyBcKVXQQAwJPC9YBdlQ
LNwpHX8okzxSaSfJRiD/8DL6z4170MjfXFOBzf/AI2KJ3JWuy/9dOv0ZJhxwSbY6gWdB0vZrjAVr
cMqfR2f1FYcQkbQNX1tJzc0glbHiz5zVqLr8/E7XDO6fUyymNR/9l8wx7ovld6AXPEcTXEjNlTjY
quIFrIcAngodS1sPaphaGFxWGuI09yRwr0h/rtZLWCPyXRvYCFHD2kATC4COj8qcxcJGW+6a0CfR
O4aSDWLTKJbTbP2a1uWJgzjZDi+9quo9ghm7qEhKOKu2ovQQncz8Vux5Qd0fIXMIAG3gRFywHr5P
x4nWusnBDGKmkcc0y1bGoqdNE+dwaF5YHYLKwtuBQ12DiTASOPj1KtkZ0OPOUYeRW79wiNeM5ptD
Es9ZiY9myg9vx5dm9BMoZmo1IBvH29+pfK6mBkne/HgheIPA2xjTWmh7gGZHz9iaBHewWJcIJNGz
QQQURfIREe5ihXHtPXicwp5nyenx5RA4UXGMTq61/QeEC4C1NufEN3L0ts119X1usIZyu5zZk+17
zCbetkzA4rT6qgffT0Ddy0lIwMVfxh4UrpOz1OXi/HQm76R/AY3RttP+b0w5lVEa0a9covwPKzaL
E5h0wcUsDIgrTr+eQnWNCUTnVyL7rp9cgYz/m6rShKbv3WWwUrUftqMkEBCZPGczDD0sRdZAvWDX
QAxd0cGealmqailIkhvDAxpkrOnLNOVLF7UYcd8LinEEwE+8puk7oXlCDxs5z1/xUb859JqRxRbu
Ql0DOzBpPdY60a6I/aYOBPyeenRmtDO2T+htK5/I6ayDN/A67VhobjcgKDIZPPSb7w/xnatHbWNH
aaoCRZUYICF0SDKAnq/G7RxMFEcYBN6Boa9dQU9i/7uCR5ugrLe2u8JPnAwAhSRkkYp+16uPYWdN
3oAOPGxkpcynlPYdmWDWYcmLkIhmo36xll/d4zeAZwf1MTqrRPfqiC0QXP/I2CHe5Ks3PPDP+DwS
N1igZ2uEd6ueG1eW5MFxgx1hHi1JmAgxgPBl60tAIm2INNRyNyN8ZGXY7VD3Xgxv3Sn8+xL2egTT
HJLb+2pdocxWTq7x+A9XdpAMY1QKuEsx5ElJY5LSRzA36O9cKlUNbkm/IxCicBUKlW5/+KL49MuO
qImx9uB3lkJa912T9YZPOI7PDf90LrHoUbnoeD/LITmvAO77QGeQ+LNocqO8RJ3v/cWvMFVy382z
2ArduOWXcohtQW7Uxr23MNwG4dl3qCIjJA9diNewJ/zhv6622gNLh9L+vuSD6SlJmlFw0Yor5UHw
JbYqxkIi1VopncDySIh25LE90C9kbOT/2cC+9VcgE3Dk9KZlAyQ8QQSNybQVpRfwAnAjyXhxOOli
KVdm0YC8Vl+VOCKEzvvG37k5K59Fc9Lyy0bGlLBZ9iaV5t98/NgTnf5xFIK3Bg32gl1rWbwlismr
qRal+APxgqFnRh2lYTmvKg398I92kZOXIhYKBcleC4qdGhvFuC1mqe1wovndsrSH7u9EwkURoyBe
mfQLjDQbK51UFTqqsErn7wdIXiSdyPXpytRDTjJ/zPX/0eJOSMaTwJH3KcqUeoN/cSLyWjHDydgo
ULm+lgJh6zmBabV24ITRqEbE39FT8PwigZnBJwW+B12Ukv13lycMY4YE+d3aykCjsz8+O3AdmCVS
EVXkmg/85Jbyt/VBSDZB5poaatF1qRdx2vIqMYmjvV1NEdLGYOzPkAVXbyYqR10klgTEECH8Juxy
DFP84NBLBr9TM3fEtj9CI+s4ymfW8HKe2uLgXY0/zGbR3AZqpGptqVWNtP10xcaeifC9fIsTKF0i
HaHKG9I4SBT+H+lKivF9WDphnQuKA6E9OWcoRR7hHzaPPwKtcFMRuSFP+G86rfUzKzlrgMpAkEd8
k/5R1h88QfGn9rMXMVLJNB6sV2xaRaA1bd3mP+9sSpQAH38XD2qEEYzrCD/QgDMgeVE0e7tHheSO
vkpbNQI8UQuq6GO/EKW+uBBOpy2tQrtk3qponFai8JioWweEGj9cSRV52V+3hRFTkKzAbAYSBkUa
eYpzkX6EFlx25CBi7T/Ne7s74hKsZNCnRnpz1Btp3ywkzd0MyIvZnUL3xfu+A1X8t0fEQhHTYGL+
cw7GWNhrLmT4PtrA4jc/xB2xOualf/Log1jVP0MCsid4EHtZhsUAQID5DvoXCgP1Ms+Puo4Ain4o
8g9JyQfFDc3AICYMJOI0I5l/ALph+U9fLuJmYa+854xzLOYm2eDc4qyFH1RZFc0YdnYWJUGgP7yR
gEobA1KUTKq5m9C2dULMNWahjl7cvpuTMVA16c6Y7Ik7rUfOsFviRjnr93GGa28Z0pPeZeUIEKqn
BITNwLVjmQSar1IuyTPP3xrSfuwgPdT3akUJpw4C73WD539HHPOKA6bs0d1DBDxrMfeFNvEaIfvl
27aWchaOCqDjqJihYdKR17vUonFpvBbe/dFYQ8I/21cTAs6pmP+N//VSjf+6oYo+U5EQSRWhmONh
zWFjoH9NGTtfQFkA0IgBq9ouIKHIClJA1uHkkq4LvTC3BSEhXstkhfbV6Uq2YpboQBGlWnTPdlr0
Vfe+kI7EJXqzh+vPincPmylcJ5HtgGOPhjRHlcKHArMs32VZUR1gRHyTYiQkwmFF3Bj/pGBIfF29
pUJ/57c12HHQ0QC4IlL6fM1ukoK595kQIZNvB+hZRlOYLhI1ZexVVg3DVH4ZyA0lfly72UMi9Lef
F4wHtNyUZsPLWAtSgUeaDch1NRfO0GahfhEbsm+M7bTQEWuNz9vq97d7m1nobzMX/6HuDkY6vbsX
tBHbFBWAF1EytBuzlubBC9kdPEPt9KENVsqISi/+kiLk907w4v8k0akf972DXTioJn7C6w6urt09
V5UpoXZqF+lbEjtGRoKHX4Mjt4zv+uiziYj2IzvkGUZXupaySuN9dvlfSEXi2RO0eeMcvAyCVeN6
j+KVWgTxaAjRcYv8PrtGHg0lDLLJBHRGjqryLc0BF5sc4PoQY4hqkTjeLnc77TZ4qn1pfVNZbZaA
thPPrhU+OFQX+0xBOACR+MMFPvnoC+4yJICB0onIKbKYlcxuWIhzHYzSi+mwImQi6TmiBw2X5nuV
C0A1Y/gD50wL5TbxrDXCBwxUPjBPALYJcBpFyjQRDXM14p+DeeswEqgDi0m4uEIX7IdOty+nmnPy
Nk2sNkiBFvZS1KZUw0uoaG8GmHYeHZ0Zxv8524U+CNiE7+eAPDfbU2FnJphfdbZBYfFa0j4NYkBY
y1Hyly09Va+/Pz3rfvmyeEQAzfM1UC41VZClTkAF4hV50G4YhRU6Y+sDZlUAtvvNiM+0OkUKh6GG
bsM4dsMTOyigVuIlLpoe8Yqo6pEzfX4t9cwL+LAjqoRocxVUhGVAS7zaPn7PcNqq0+0ggd+ouG6t
MmJRVgV42inOhiQL1pOwIEZzh8P/ZBOqisWPBWjfUTsJj8HfMOt3W6tfrIocyjR2hfXIUR405116
i0tFE13Yat1LQw0TJCFWoF8wqEuSLe5585M3s6NKy4tpSrLBcC3ThonGvcKL1shhoj/7e7XXJruM
yon5gjuHhdHe7BIPICAHYypS+fwdqrp9C7lVFIR2a1S1So3efjqU9UiejUj92jsbR9Ytf2DM7Ozj
3tTXwICSheIz2p+QnyQJbPf67ea2tqCmm3gYiWGHdX2ULoAp7lHC0gtuiQmDNnDZAQfK1LaNBhIv
lICadKmn4onhRYMOrp/3UrPFX2aIT/2gmF47sInlfs41gEJ09ErKyJpSFCPEa8dQETiJwMrgqpU9
MDCZHzaxFrL8hh5nEYZAtIwzTVaWTxk2wiu/QI0FOBECaI8TUTggNSM8C+8y5D6kKVpurpPlSIgi
9BIiqWt8FVmc9rozitZFR5xYxPhuTtyHLN4M3rZXnMXin80Oh9ViiB49o2hEawu5gr5ssywsa7ch
3eDev1DnSfMTO8Rd0wIhFB4irr+f1emQIajw8UY4nylbPzuYl6FvEMLBKhmSElfcgHL7q13qf2dD
L7kwXz06zCVXBbGIWW3iWfRRUhw0URhg1sYLbfEov946jWuWnaxw2sfiVg2NlvRxyfFCERWKq5Pg
wfRBE0+LZJ/SoXsqG483k32ZZzhFkGcFZEw1/QsiW7DmQxhfEAHXv3nHcpn+lyD8DLpdfKsFoqJJ
dNm7Hi2i2qb29IQs1GYB9tb5WYN4BzKIHVgpIJOfAB46ByILOe3Di7+6QAhPgnGtmvvw7PU/AV3V
ZiDaZU3xu+orK1Du346xxrGExxp2FxMZNj64BhgZdNCZ4Q5Kf6xVjYdMFs/L16Nh7+y50u8w54gr
EUp9dEjHghWlzFmuZESJB3d9DLk11lCt7QzAtyhyjAxZf21BgvH1VowvIR6Q0cVLEqspeq+I3fuY
L5Phv9haxw1h2JlKoxL6t0xOStqzwAOblfJETC9ufV6e3ZRFENjO2CjJ+cwIm+MSuENxnxzfDWY0
G1KhJa4RqtWV738+vKmH3mirgpZcY+XKxcjqye3Nh3Q3kEfEBGhE4ic1OXV3+DIxlMdJ3j8VSDb1
1H7tnTGxTi3xM8kyH/b9q+BuXdvh6P93DQCFtD/XV9zA8Xz2Fg6uzrlXQYeHncGu84hz0S2nWbK+
b4tE8nLloAKWTalxtqh3LRdvGlmpLG+lNl9JLpvvpsJqx5elFUPVfILT88aYla1qTIzWcfyLRrnU
gYYqgO8E8JTNIkI38r4XLmcecKDCf+CO7FrqkjvHgv45mcV/pyl1Prvpi8AVAfU5i+GC8GEzgE3w
V3geCveGm3mmuMNV1BCcmT6WczNofxKjS1PdXH7lmDJOKFecMysGUzvcj9lBw/A/0x81wuDXGvYu
vbTxINNmwoNaumcTfcm+UtzhlYVBUlg1Prbwypt0772VPTGsu4idvyQMrS0eYE8sVE+H2ecVxsYD
kPWnAsKy7QdbMJfQARELVfgKYMJdMwW9SKM/pwahlnPzOoJGIqyt+WsNairaVH/uTS8vXLYqOEPP
7JJnh3jnOCfKu4/P4nvbHn/OiQB9UzbQ7dfZzEVsymswdgCvW5oVZXtBLvIFWBFEkPWfgrtzq7Lv
ujMuWmyyO1naX94cxmxRY1ytqZoPxs603sNhMOYnX/INwWSyfJkIj1zJvmEOBZYqHtLL4I2IXijb
YYiQWSe+3XorhUjSb8ScLuTQdIOL74Baf1rkkGV608yHn3SeF/PK96TTGXNv8wP6sFCFKBDe67im
QG5wzR4J5cTOdnhNwj7IbLEWKaN53bdMTQnN/GR8n8revjRLSAjLFmKBUPU9Gz65xTultA+TG4c9
ktIkZ/QVPcwZFTZMMS9tRw+n3irSEfMfwEiIsVywa61Fq3hFKE9SaJl6CMjXQRT/1eAYNhZxzjNR
gK6FDai9CLA4TTaTql+eNZRgT8f9qfFVWVNvV+tbkY+Oa57UDIEN87h9tCJjP3aCgeElwL0qe4Lo
jDqjXB23eFk7D5P/FRep63RlPMjKUHQGNSU7SDzqNHEJmnvduOSd+SK8GAUOtehdXi33ype16mF3
IinHEJmRps2Fib96yZRKJShunOyf6kmFeGQBj/6mkaxOURfo4nATDsVH1z4xM7MqpMo4d1DL1b3X
HbKI90u2cMO32GOMGanaMcax9LO1b46AFQI2kta+JbxsORYqz/NH6Bwcq85tf0K0mKZg0jLsqE04
FePg2g5HhhrO7wZjOz2RUc+WyJtpTk57Foejg7IIEnrqeexUKShmOB/oEU25KLf5S68VMYld4Fxk
FZp3iiiR38qqnI5kmD7+Fle/SfPHPsOzdqmGnMGtGxoUePoIzzQvcTYPZ58CMcFzhomBvxJIPkqg
UhzsKVPso0YR5Jte2nEnmxhN41dTn2adZ6pgIuYb7SmdnRJv+CRUiTxCPpds53CYo31KryStz/QH
Y2nLQr8me7zRbuDexG6pqp8IB1JTVDeafjx3zVpeposWM1AebPgKfWx67J2rVXQqeySldWSl16g9
2u/UlbApTIx8u/RIaF+xzcEHcJ3G6GLDo55/JPMQtnaxVpAoDwokTdV4tOTv3XiUVv48xQnS97vz
EiXqO1D2ULtHdFr0r3p5qd+YSaD8b1Mz9NGKXP3aO8vVe9L07a9sYE2MoL+qPTUxIIHWi8sUB9GH
5C/MU4Tf0F/SPXbSM8lbNY4DbkNr6GlDldLQhsTx2JLIne3maG+hnqyLmpAy0z/EgAu7jx3T3cJx
cCbYZh81H1ZF2AIPdVQkmIzunNskG3mfbOFCUtZOSC+YMWQ9RpDAn+CTw2XfIuGho21y8cFYcoTA
SkDv3lPxeRogkKSliNgjwDOq3AutVpH1oaAUof3Y3hltqeHcvg9Gd+X5HPcyVU2kqK9PcAJUoyIT
5fmbo+kxR6YFEM/wYHiERF5ogGHDuMKhYOx0tqZh6+rIYCOOxq95zSWd1Bw/gZ/E4pgdEhv6pIEn
08fboCut/80cZ+gAQKoa9hQaASIupytkOs3LSynUWYenYnhyhWDUT3oxAEZAPmflnG4nT0xGAkl8
ESek1nc188EItcfY6EdB0GXTWT1G6tAJvWOVYgGDjiZH0N4E5VkTIa7VAzy0EUB0qNShfYJDus1V
RUgx8bcxpG7kBr1qskZ1Sy4GjADlCMwmGG41VhsHVm06zCsEPKLGjTNEr8kY/4+Y/Gj3Xq4C9IDJ
AZc1Hn4Rp/vCbsZpZhGgJMKY6JwX5MRhRrKcOxNmhPi8S7go4t2wQerJBJLuX4QIQEChmZARePJF
yGP968t+4nyp98FN/qf897OF7CqaJqtbviHhXx+B1GtwaATyF4skWO+nf5MRztWlChuFeUa8nXYZ
2qKgkHF3LK0NrgbvKJ7J6SCtHKLiZjMCoHg52Cy/3mTHM/+pCJcxNJKRQrmBFrzueLvJx1wlWJRa
alBEx2RKzLsfHzWmD6cCRewk12NFyRFiFthsmYXGi5GAFsz2kaDkC/3VNAuD7QFf5t1GEgJUNTqX
5xkEAQgFhcIl7a1WVI0TvflBcrKnKslmJX0JTY2oG326LU5BUVacwsaRpqBfDC6UThSk1xF5r1v6
mGP4cUE7sF84Hcp01xkx4LGMd5+z6VjSCgQKg/wspdbzXvEHw3gJRdQKdEr5ABdKWElmlXmEhW79
u+929BHgaXHNo5JwfP66FpN8N2Gh3qj8/+dkNatYI8Gpqqw3MOquW7/ZzwKMWVL0u/YfAwY9OdF6
RmbQks4qDPnoJbJM6HrpOuw7RRqksxgoE8EFxwIJUsIlRd94KINaRYH7CIpaP+m5wNrlGX5yM/Lc
yeJOjTG6aOzjs7WOIej0uzmHUzh4g2hrZvYJx5kdgqksZ8Px7MwHLfLKWDXpTV+4V5sbQvp7LQb4
6rEOfruOo6Fq6G5AfGiTLBVM6E10mIdmAzifg00vA6qPzAfRYwNliXox7xul6uA4xp5TK1/UzMJ9
/HRIdE8gqieus0zjTX7HDY6/lsOtVrkGjAR/8kaQtWw2rajJuEqSGhe0rWSgDvXHL8EvMa+/ok0Y
xI4ogkdLtMwBLODwQU74x+rum+zhZMDKlkdJwhDoMkL2lE4ARilx9Kw5KU7pGq8r/2JfbZRbur81
nH+DKFwubcDMV4iahjyDOnFS4eLnI4CTRCAT3oat3ZfjxeA6LbbLwDJrttvjPQsy2ZqAtojQCm+H
4oafhLuUPed7YdroxY88N3DqdlPvsQa65bzxVBGv50o6WgJZwuYYMGtKIh1q2w7h6bMUP7R0t3F5
egU/Gd6E1+i2gOI9plUksYojxw+m+6FT26KkdCh63vTXsioFoD2r2dXoh8sp5UHwxDRMphTgeThq
0JBePApfwZBLmM8hHahmH0vjdElC+733d0D/Rn8cl5sa2tlXoUPrZKLWVC5T5dvj4jJKnHua5uXb
hgv3rE6rJX2+cLzGuzX0Gv+05SeIwuNRHic42SVafmNEs9YzQ+2qfNyDDkkYwl2ZLr1u75bewK6W
DIwgTRZuKLxgB5K96a7BXK3Q0jGnRAlimUb2qumD5wIY5lZ7MW/+VV4eAN4WzDAiu9eWiAXHuB6l
SPksQoMKVSw8DIWndDZVebGhloPTKqKTvyvXW0oVd4uNWCk/gxtK8avuK1+B0mSj2hEyPuB/RTCB
QFwROnRhc+MreaDpSPMs8VF6PdhM0ajgPEkM1jKz5NSMzfMaGB+7C5YMXfjYhW6DnFmyh31QXtfB
uLxGVLWaPTXDEimf241wLmcJ8D7BADrkPe/JMGNRnSriSazmxzKkXCNFVeDQwRlj+a7+hros6PTP
yaALwx/ZHygt7FM+0bPNUQLdCbA/W7kK9Jsqt3bOjftC2KDl5FSBG/ptHlUARTDyXWIVOPKil7lN
stVb3o93SYFrycxOC1uOQjkvlHocI+UJb6CD7RzkWCtpaxnQNdviP6kb+WE7mYs/ZiJNUgTD/NoI
iKLOn+F2IA1XNXFCrOVf8cf5IHKAwuNLhS0TSqA0J+SGftWWLNJbaOStpqQER2rTUwiehsHEmq+Q
cui3BPUOqs/B/35llUrZwVl2d7PIyH10w/dmQVlQ9WkdekKfEchHlip6pKT+BftGQGXwFEGv34C1
uFaNOTfkknDpzXXA8Lr1fKjFUK6STlrimk/5R6JoUijKTlbcTqzQ8aUfr+oPzlOLzLMr5igUlSDc
PU7mNGx9lmA/tDBp0IqJo4Hcy+wNZkM5lqW4yFwXwl9p/ict26IvMghk2m4hiSYEcpqo7Dp7jbPe
rYX+YWZKiD5t+KCo3QW939qf6XIWjKofftg1GYDDhcwUJglhvCcLv9ns7WeAJqf5Fc8IlJTWmU4P
QZ3r43HQj9GMevVzeY7DW+lDbpSbdZ6G9WNvzkT1Vx5pDfjqi9a/L7pR/x1x/kc73iLWYTOuTcMn
q9zhiOl6/N4XlfCN9iZjtGOGyZbC1t9Og5gWTOCoslGlqynWX9sENhSxOyr471Q6RsR35aU6ztcx
HGzSEasDHj3vBIO6hgtsLjqmdQuzXGEJAiXnrLWq3sMx/irMCHaHiZzsCHQEC703ONfgev7Iw/Bp
5D6j7bUlvjI4KR0QpZjE38EsFZCMjlsP8PGO7w6jI1dBQZrP+3v3b7s0Oxz4TstbvItaMl2POkWf
j8lGiCxGzud6CyHkOnHCCBaFF6BrU2y3d6UOh+O7LgItOH+jFCTsKzK9Wge5fPptkd0wFHn/MwmQ
pn9YiXayoZ/ZbM/1KO+FvM9KTM3ZAbE2WoPvHeCR7I89my+sE+X82DABjt5rwSHw6roXsksK/PeZ
uIvnzt4S8Gu22U5B/pczI5I9nhOZ9DQ+L+laFt824EFhcSlq7B5RIwhE3T2VmQUNJ0c+ao4B+G+k
2Gdm2fwlRQel81PctaaPaAE7+TzenaT4sWY7dOBy6TZPKMBlEK9gnr19PUP1vkn4aPh8i1UAmzwr
sdizvjp9wRqYM/OsfDyVSg79xvQCez6FFxD/SDgRg5xNFoybwWQicbVnkxadLBeG7sMIzDVweBEg
/UMiDzf0vA39nLm39PIg2ex/bmm53aJaUcWDc3z9elwpBGxmydQ92h3msptc1NBFYVN9VaEFvJan
CA6V03FUZgcH4tj1wzoKVQ24k7cFqbxo6snM33AeGD2XEIFzlqwXGRfGveckrAotFy/j7Tkcu3M7
LPt8I/qTZG+D7d7GYriDfJ2DOvRYFyAFRuJRjyfV+UufdPTNJI/fHLLHZqhfgjfxD35xUchDXaiC
U89iG+q3FctG2pNFcfZiQmgLnOoBTIoupRXdnYUblC2AJIKGaGnWSlLGkCIlmvhgFeTDYxJXRC7l
mA/Yuii1RWXz9Grt2pNYC2457tez2PA0jU2ZxRt6qN6/iRSSuvGiMpvrL26N3/PckHrlrroZSQ4u
oh8A0yf2VGcZBDgw8ymFLy7DRsxDnm7qIFg858IA+wgds0uQC1k0cwSxx2nEjojAG2Bl1anMJ0aY
kkc46QQgdc9SuW/Hgj71qf6Km32q6qJ3FfXqaWE1PiahWpqaRFdRfVwGcNYrzGiMLZ9VZ4lEaERy
6fKqgf1R1VSY2I7hfGIXGLMy/H9WUyBfd+y/akAIS/VU+hNx3GP6On1sHzLANaY/WuXoa9A72m0F
q9fG4+bmwDiHB1jwpSmFdVnWMmdKHO6/IUfizVc/668795jNGuy2cVIdH2btAJqPLMAt+R2RosRi
y/xWu04N2mqnT9UPZ4r/+1Rs6nUBv5egWzMQrV2Ld+RHc/PhLd+b813qKqqqQocdp3yPWi2FjnL5
uMFIVBSs3Ec/omhiQzwuAEZrpPda8/FjHb6CMvvNdgRhofziCUtWAitCW0ri0xBUzya3UJZQlC2W
4r5oaZmHCA6dymccgg2+idf+bQXokKuNzFzBq8gcV4xIxavoyj4RQQLL8wYlMhMk5f0PeDi7mv2d
uNOKMVsTsDTZ4P6Eelg87Z7WwIkzpgIGBQCNVh3hErG7M9FafytBbOfnqTfThnSDSGiUx3j7nvki
wpi1RGStJv4wunXrrtw+vgqxDv88k+lxgovBnWON1wJSbZDV7BwjHZoYcvB0O+3//EvwikZMXqGx
xsnEvzTPP3b9g5nsMTYtQbrScjlMjnVcv3mAGidpz54eMi/Jg9PVsoEqp2/hCcTW3lxMva5a/G39
SwyKkGDKgdOrR+GspMrVr/KH1pt4wFyJRK5HcOLyvqT+VY5kgdMpVM4u93JqhkA1fSqEHP9OxLHA
l3Qb6zTHYHTZ5ppNQFHghG5T1wBHDJ3vHYHF81tjHpaosGS/+MpSK3Q9bBD0HeW5JuM/+GDMbzvN
SFU6gBCPgA+eC2R7zaSIH4QGNw+b1VAMYFbk5pvhwOszFh62E98JibUO/aJMEnLWzVKeGBVNYnaE
3xQHvHugOtr8W0hKxYP/PhHAEWTCtZlxSZRgrVFNxb/B0UZbEASYng9kmugelQJHbdWjFiPzSmat
o8kXHASeC08rWehoi3Rm6i7nKutAoxTYsNlC4DLSbw5mt/gMIEtm1P4FlJlZRtwBHuB7X/ZWXV0C
tXEJ3OaTdVkfDgfmrWamBBEGKPcNSgBJrKVmp2bQ4w49LkX/5mCa1StTuabQz+1z69KZC9/AhNbm
w286d3rl8hNUrswV8KRoJ9DG57/IepybUs0Q89WHg0nO+v0ZnJKw4EGKvG5R2YTNiVVtCsb9cU80
WxwnWrOWstBJoHuOxESrSVdndHgZsl+Q6Ddae5SaTxcDYFn9pS1Q8JrzHwyP0myUD/LCoQUHYg8S
58FB4Pl8m7BNLlbAzujFkNsdK3HofgP+uEg3l3g5SztOg1YOwR4I1qszaZLs0v51ItLqcX0BQtPn
WTfOWWje1MpPR5JhtFW7CZiPaWDs2ln8hhxgKk71M33HQMMaM4zOHmrMquLReZubKWot8gX4OATm
vRvAKhhorXLTRLloqI0woJbTLzvgvDWDxHx090DchRKSH7aA01+oKtTz9BvcfSPAAOjw4bzBFF3L
Et7kWecVdLJBGLHYQN+iWhB546aEXgMbqOsSs9AobtWcwIlMSJRW0EkpKsVAWJCIG6xXGfqjX333
+2qUJ3zN/pdfqV51ufswKYKD7fqGjFSBAXLiX5Qp9aVMV4OlX46UsXoduwqe2K8A4T+X8cx+zi6n
+soDAhTRZjchidthBM+VV/tCwLK+UwM8W5mqKsnAch7tX2e5ItiJ8tuHxCkt8ZMw8Owe4F+TaKqq
u+mlJKCB5PgLnhVBU8mdBJ/JaaqOpmGRXBsZeoQAZ3RzxYYF2WpIF6HF70qB0YC4YDzdrC5fZZQh
agoQ5rBLhKlpQmLsGwCi0min88EygXsobFGUsxgqaBMZTJUoBPLR6T0K6pv6IKEOWLPHLXj0VNUr
F6rH7QARxsPhM7NuVvstElOr7c+QyMigQO/FfwH/LBygRufO2p8ryTbCcL/Br6C/ghNVITxY11u+
AHTcAo6o0aJcIqLEr9Qz4E+1Qw8ZQ35XZKeIezT4a9DfG+nDxsYkU7xRDb8/vQLS0HE16bNoS/Z9
s518lOfvHLU42hJb40WJm1VmAuwkFTl/Uf5FTA7BjFeLAdEFYVUf32Kro7gTq7z7w9QN3MGTCF5Y
+pwWzhKWBeG01zeytuJLcFcjCAQhBTNdjxHvgtfm1rLbMaUnubSEKAQFFZZBM1xvKgHrmRkC4sEp
wJs28PAR8riXUVDRZmbt5Bx/D7i19YPUiOukFkRuZqwjlPrrsuMlCOe8iURMwi9NP90fZYHCbp9J
6zLVRLZ5lgFDTL0KAiLZ8DMVLLPiMGSdXJ2vSy3Mwjl4kt1g1XyZ9s14Vfm+kvCAstADS5NGM2SI
/gA1nY0DXgQaPjZwdOG8qPNVf+8L5sZ2lLGfGkBgky3zYlfwyAlAUFSVJxbghuBj5RvVneMHxT6S
H/aYDtGcM1xjxgE8LRCVsbI96bqSnCBPcq5+sKxmsc7SSRCBy8guGoQOeHTGEBpeK9nt+jHfZ809
pfL8+aeTzNHCp6hWs9BG5bgUj36IbziTKDJ88bTV4H/j1X9bplJ0YookIGHvI2qFg+U4zYF6VMEq
jboVPQVimAyUuIF9P97WLNF9YIJCytzGQm7wJmCkrSkJTAW688ulxykwoABCyZ2VM7ptEYT4w7uk
ukAAL6OmDFtMt0dLeFq8Ybpp1XNEMJ+NEA9KeRJlmiLL9DS4g2wgXpuFCKU6UEOnNEyTlKp9DEI+
x7jSqoOdgFkmtKshSXazMM421rRLOYe15jNeSqoTxsvW3nkUfWKE+UYZEze3sdos+qAk4ajnz2R/
CYGXKI1e+Oe4q6Day52fVBCXOCuPbIYyge1BJoQ2/HKc6pmxtXPjZ6U/awvuT5PaEWmFde35s7ES
YpTTVCgq9PA51co3rNag4G3YPiMv1wl0p9qXVGNtTsqW1TWiaIc4q3Q6RCYMOGCphUcmGTy7gAce
P9+nWCaaZ8rwuts0dZPlR7Zlf+wPApj9R+IZhProDNrxMYXiA1AbRuioeDMRvYv1kPxv4/UADCUF
y5U1q3TeSGEwOXJ1Dk6QLTj3hAvCknW5Y0OK9a17FDs/8yppxEeXv7ea14REa+gNOHiTZA+EY82n
H2tpD5FQU24Lv0skiGmSiXv1G07hfePNodHUBFNiEw0v6JnkiJcvcBUkqTnBDeN4luMvhbpLcVZw
BvWbBzA7NEBUOezqlpb1AGFtPxi4/tZaJ1ex9eJoE9rquU9obXZfodq/Jrww/pptipqyG0QgO7an
NP/upRXX2NUm6F91hZzTG8XVARFftc6TzaAhiMNt1csAnDBjheRmIoMkkXrl097KrwzIEyF+7q4m
L2CEnSDxAnJQKK9RhBjJ5K2FDSBTcvRf+6xtBBgxxyHtD5OOM3gJoCIZNnJb8pgFPaykDWIwq7y9
qICvNwjygkBjJW4k6iIYK6ogHPkrfHEfAOzYtZiN29bPDK5irelABi3ApkcYAXdFjrCzVooQLxpS
fxZtpLPGR6G2J5eRqoF0riBuQn4qCT0zjo9NU8aW90eIwilKi4vy4eUXWivdObNw+OZHWfXE/O46
2RhIrasPlYymY9mf6l+FU2bCbzgKcfIE9WgvB1TmO6GcSCi7Q06gF7925TgU/dTv88cD1rHewXmr
mgeeA0dp9Xlrloe/b+PmCsv3j7NIE1l3EMMcAUkEAnkT5qZ0NA+tjC5rAkz6UlZdzNryGLexveHd
AFSlI5mBHpLne7VFq6KSktF+GVIT7V1VIKDYlz1tvZwOMoSX1J9n2IowakCv6uyFvHSE/X3yxHij
SYLxTtk4rXdQWWnuCzFIWtIeFETgiu/8s5xQppGH+PhuFoopaHrKrlU7XzqQoBuLumrVmRZ+iUQd
xVRfsl0CfYpLgGHbj3XgxEm+OANgnPtfjx49EDHSTVZE73ODAD/ar9sm4U0c8DeZ5fTZ3ax7njfG
PszqyVoE7B9be96duRMLfy9G0h6VoODZkI6GjffSRcPfaZWcqZgbaGrkrSvuuBJsAOhlhEVJ3NH+
stcN6SW2qnDtqp8B9kfrS1mrRFYfJT/H6PRPgJ+/GUwP7Tr8qYfFLGDNy6GjQJ28eQ7RYi8v1C1v
OgE3x5xeTwX9fDi4iQQJdBvKlFaBFsVuYNXR9Ab+jAFJIBKFZxmfXsIUJ2rTLTXtTI7+mGwMsu59
PitjvbMzMv98Bu3ksaBZTG11ZbK/O0JEazDneV4yFgG3+7A2vRdDS1vPUHrzP44zFtqkFjsfbp71
avYkHk/mDa649DjeosLyLhzBmL0RGoRF5DCyW793tJAX1EjG360NOFLkYpYobO01ijPeknbEFnfq
dsLp53WD3gdWfq6mooI/1uISXa2e1F8k/tFa7KaTSu15+oTPotiYyZ0Jhman/p4Xy3B+Ld8tQy8A
UH17fKN17T+PEk80rMRuuRunVnk4w5vlS0H3gNLxH0zEmhXoMeIj67ziS9P4vKx8sNuRP+7yRUaR
JkmIU4HY3IlJY7oMPcWcRfekvwRFJ2FIMPgfytuvFmscBTVRFvmzdMaSevCOswik9X0QBAZhRAoU
iOlVQ4AjBwIdMVprU96KqA6OxtNHpptoKa0fIbYLMGnPqjvhwkKmYDSYkG5LV2uNXV6k1aSZVPhP
eKLKFmLUbOA5LQ/btIi9Qrgs/L6R7qMGk67i6ssw7aFLlESIKd+F8P1xLNyaCleEC/0QRcXMgiHt
ccMYfjXZRGSOz6lxJpKqOTrAnb/wpVvTvmoxiCvxHwJeSFt7uAq+Z/3zQ0N4XfQUDdBNrZ319qpU
Mxh9md9EYInY3rd2iiA/S9gz2kXb+p9htC/xgI5ATMf8itb9ZoRJFwh0Kelw2Lk44BwF1f4uaiRP
k4yH0Ilq505645Wk7FYiobE9/gSYjp2Wb1kgZBo108CWXNu99Cx+m5FGS9Go/jCsGGccH9S87p7F
BXvKinh+LaM94b1PYee2KaZjKUjI+7pNRAWxPymwKLcbPjl+q1ltzMOeyvFzkRQ/rlicB/h20owA
EdJvWQKOo3HVjyBzV6qsJbOuW8DXHrXr4+Axzo1hJnm/SVpW+vumc+u8NAmRosLNTM5Tpn4iUL3v
7Nem8W8TPb18fdT17OazQwbXctMtCGUBXEP2VxVDCmp3XTG82uUL69WA2P9JWE/fDxd3Jji/CWs7
rVwi5brNMhxgDMXPxRB6cNEHjLN1jZSKym2pVIMH3At9g1mIZzP8cXbpAgDOjuMnv/y+WHPh22pT
EXu17ZWym429wEs0WK04vdANtx5Duc8/zkW26qMjyI1pj8f+Z5XvPYF1fmZT+NdJ7T/Pav7OBrmH
B5KUekZWZZQtyshs8UlYeD9x/pRpWwI8S2nFCqAGcCU1ven7Jo4Mq/QLO5wZCSy+bnvLyl/gjzdU
GOiKSQSEfU8ykzMibei041QXEwlpajdSxYc+aehPd+YNN1EX2LBoj3oBkqZEahNvemcxHXVlFBxN
a3pq0qC+DjSjkJk0g1vgRVNIREpdosL/hhRuoHBX7tDGQGp1DrphyXnXvcri8eRiZ821Qpe7sCY4
is/dZ7vODPyKc5ahdNuDJYqivgd7cHC9bG8aONHsXConeGx3SA+9hrm3YyiL8TYXHW6WOvwg7bbF
HXL3541FsLnHjGLG2zq101CjnqjUGN2x/9y1Hqlux/oidaiYj9ymIdvZ7WtGh80vSHpoFCjLcxS1
shW35Wyf88qmC6NX1G8iQmQdaMVNssNWAM39iUj2psFB1rp8jmi0WcCYQRsG1OJQc9jBB8kS5JKe
N3TitvnzQ1cYCqwlAsCdgTAp0p8+UV9/NPjUTt8d31RnfP+5o40GNDeOYRi8OjsdfJmQQ8OK9p9x
4HPrRFJXDqDJ0bQpdiZI98F72g7/FSqG5If/qwFOu7cGQhiiYiLGEfmozziibEd8U+qhDuFWhHR/
DEEGfTqeiOXdGGveJbCORRhh2aKAZWPd1yuMPISVzfIbcNimBfOaN6MD+twsywZTkQMXq5+pEafM
GJ1dZkVLxnQpgbJdPXiIMGurUoxmaPxh8EqkC1VdHfa1xrjJnHjsGmFhUhFV5NykZ1b7XHGHDWif
6vOXYG8EvcKnHnnP1omhc36l4Zy5LUqA1YKfOBC9a/OYJE2U8EApGdcyPFJYnIn6Ipu0JcKr+rg5
ZnBne3D8lEFkC+VATzLc9503jW+V31vD3jf5ZZscFxfbX6Ht287t0/hykWS3hH2fwAcrurcCUIqm
i/ecgoiBa4rs5tAsGQUSz//+en2wgeyHs/yP4HnyVnLvh7zUJ5OdJBYM91om5H/Ac/tK/eY9KI72
NaGz1kU6nKo/YgUyElBY0xRsS83LRZ9ORg5YTexNbOL5GO/Q2VwSk81wyVjzAn6wv+jU0kZ3FkI7
e2iG3Fc7cgD4lKB3PkowRXpRA9Ba0c+DsGvbwtbH9qBTr1sRYOvuHC6GyCYDVX24DPNelcPinAfK
XPezYrbNaSzgOh3NBxdr+/Ei1pyHxXNdnyhZZEyzIuUhRUVDJs9bQWi9euTtBpMYxDdG1e3l2vqb
gM5e+e8twEH8HnUlA90fhX7T2zyEtva8fwvuueD2i4EYKnAokmq0OcfGYPl6uif3bMbfTR+LcD8v
gpJ3V2IUPECXhpmj/LcKS1O1e04M1bjO/97chzNDdeDNSomU3eZWCU+LNIaIFGJz9HonNKdFl4aF
azs7TY+Q7+4l1OKkhmzilZdaRHTOdlat8eahBwBC/Y7e2q4Gh+tzXDEaXYg8iJkTOn6c5F/jXnJR
PVHWEPJ7U0nRTYWcNr16uFKLzAXC5wSpV4DM1kf46Y7xHyDAj9fzPHkRFCjtpeKbKOXhtwIRjzvJ
jQviJUi0jBP9NekVV56XJ6kh06qgejgYu51BeFOlKXP9nBhvMwX1uRov3xPgkJekHGySK8jQBNiS
JaSuOjClc6PerKZrhJ/Ehfgncc7G/19f2/epMBVzT+8sQkD5u+yqVsZuQNwPDtL+7d1iCpmDJLTY
juUJ51jFB+yss91us0lgZ/ph8ySpfkEcY8XZXK5VlPIA1ZQFdOsphacbYaGnYwZAqQlfNeFRsDFP
VzoG13Ng99+yHlc5IX2PjnmK42JxLLk8AFc0Sj0dvNTTSxEUsG9mHyluoXhouS2WHnaf7YXsQXyo
nu7TvbXTjojPzi+GOoSGzGCNSOLUSYuFIBfrflIFmRFBz+Ib2HRCXk6IGpXzcFX74AlaO3Vmqcx0
/LeYMXwA8o7rUo4IZkXQFo2+qbMIPVA9HZ8jvjMZ2oFD20bRKKgq9GkWzb6IU3sezzREZo41OFvF
qnpDbqOMM3EnWESiyeKQLifE48Jp4GCuiQoRnmO14KUbXGaiwnhC7FKRDEGVAhqbpLG6+oaOh8In
OIAkQ/sQcK/9IscROBJonrXUPXay9RG2p6q46ljE5oHiMpFqtOam8AwhTkU8FXC4WIa+kzWGk8/9
PylFeHI3CWTXfRm+PrTjvoz9L46yq8iz4G9AFetogMPAPyrVS8//dnTp7pAwJUesDuxyVjAz2iV9
SqcnlaBuZjjSSt/tHvW/zBsq/ExjUZLM64spwIr3m29Owb6rQBhu8lkpEBF9dit9oCraJmfJby3z
xo7LKEhI/qSXPYIKWvaRFxIPIDdPRP4lixqYMTQ2df6oBjm83Jl5mg/Dhvjg3XmCQC/X5r8X3E20
Zy1wnAH30VTDa74BRN1OV7hXaQ2jkCMIsjlfE6hLkd/eRpG8/cNNLLnSC2V6DlWO+4EUt7eSq9L6
RL1mjvIo/9ucuwuz6SbGXxj23C3uVhG3lRGCrRFxBSjt5L36nAhlqwI3mnI/jW5ewdKaEKdVTsVM
hIIHKxAb95vsuxOLrFaJGAyQJx7+D5GsXcp+nwBSfDmsPbFaG2H79miwoeJenRxuhOOmnGnLxadb
WzshAhVXD5CBilhRVoF58K+LYv6CvqBgwhExy7pBhwW1sM1TvPqFYGLgJZ2h+oyFYRzAri5reQy4
Nou7FK2ymSPD52+59IeURXIdNXDVD8NZpTAC48Q69WW47ItW4lCZo4heEEz4R26jYLkPGcTR58Dl
BVhuAPqPk/TTCGVqUGMygp/XqCkdceSxsAyejiIa6PPzS4mLhWBdhdEvzuI2boe+XZb+xKLHkrTI
NNrznqMSVUDAvEzIL6HTqZymzdYFz6g17qKf+i6Jwhgn2yF1HF99NIIFpHFi5IEzdDFADouOPCnz
kji2QwIVGU2MGEz6Mmcztdfw2FpA+xm7h7cOOxa62l03kgAw/SQE000s+SnE8CnNJB9dXqnHMctb
yMkQj3zF//NSXPXSFgC1knpfwQa5phAGHaFVw6SgzJi8qrDbW1unKAa3FVZREN5yfVDe4bty2Su1
jmAIRs0wwJHcrHqZyL8bDxrqDv9xFXXxL8RpTPbE/GOBQZamoYMGHMDkUfWulxSPcPyHJEY43gFF
Nq7Nk0EgJsegUsee61PKyG2QdByMqAksrgL8d9KF2mIEWN0zaYO8kKPsBYp7MyvblplsDN25w86K
GLHi90BqpfDEb0ftnXCN0yWrL7GpNTpgsVrr6MKOV79UNq8olORM7LDrau7xzTKVM0SVyZJilB51
b0zV6pVPTZrIqrW2SZQEvUv91hzmG9EpaMYn2yALCbZVCHJRs1TFGK7TltbWjzDUsrAFAuoQnQTV
HUPQqoE2EYzljbKYKH6xVSHkAzPcpLn9cQujrrU7yRoFWJr/8h3r5uN6bJ6YRtXDnDIPU94f4kVz
cv5Cr9LKgnQNe3b9JnF7gGrTX6dLTS525QlYclbwf4JMfVl1cNY/Is3wGkXz88dnWReJyVBn4P5U
cDsla0a45pkKJKSfygFQP01RsgXhY3R7W8YANzrQjkFZlJWXQG00ybs1QImpSKiUqSYjAdvTsMat
avKkU5/NJ4ENW8wDfsMNuJZKAOnGL/b4Cz4CQCLAsl9EBMAmCuU9oTDxdT6kQ2BB6EicUUmK6GrL
Hcozru1wzdD3VthHTxtVb4rxIF1A7pF1+UpvwAPdcHtZFAN4OegVLYikkoybdd3fJGE9543uGkHL
0x93pSgnx1exGSLuLh/bhPJI3yDYHaTYXLakUlcWBpYb5PQcFbe0wTe8SJT7mN1txzKV7jxDYcHJ
tbKGL2fkijW50ZnOBLuiIOcE/EdvRWtXJ1anSbhobf7ihfOXqtkMqkxkaq/iOX95D3eWfx8orakK
BzHB6qYA377RjZzea0WJck4P2oWj4Nyg5j2U2QX08t+mpmFM0XH9nNmuZV7odSTkQ3e7S+rWPK64
e+JrPYzOKI8I2t3R0I/MxKyYndQErHf2wXwPZLNW+gBrTDZ7DytrkbMhcWcMkd//w7uuO47qmWVQ
8I04dpjreeW75EJWf21RRXxK//MzKkVL3HS7o85GCECfIwYQZ/Pg81342qctc+4YHlxxNXyB9UH3
ksVYtaUaSQ363DGjUxtvVIVjoMAuYq4cURPx3jkq/IV8bNk0lVJRtK0un89uZ/9996QZRgv+6r+g
vdWEgxdO3zLOQIZSYoyST1z75LenCF/8zX8sAeb6fZQrfqwUd1iv+Q6OBswGM5cZxCbMIwnYa1Ck
h6/0Q9LQt3JouMYsgJkL+fveiH4YNPXIRN5c0sJKMTSJOdYB67TfDCVh0QpORi8Xh8NMC5y6H1iT
Prs9Z+r+c4swzMyQXa0lExg+xktetEdUqPNZGyMFCgBxHm6oXY7zu7OjBWyfnpZqDkBUObtKKcAz
42Kw4UX52atpGt9NsL6o0Xk/djyd5zC26fuV68aaVNC9vUSKOP3fBTqP8K3ZLtF8d+bSw5GMLIxm
Z15tmon4iWrRN5Cza8XJOQFVmyigLyRVJAyc5OXW2qXL9nDlWHLd0W3d1ZNqr+f8ckv6jAcfkSAO
BFLHILJCJeTj+IwwAbEgNmdf1Eo14+ifpOdTEgDTudNvoiCjaPSJYzmvPM5bCkwqEO/1YsZt4HkJ
6w1IyKpw1EbEuPfol2vmcAndUeKw7V8sdlJS/g5k8BTOI2jZTNchcyLb1O/b1MBcznlmQjOUOn1N
gbTK/XuAaPP4+AIKb7GJE+KRKlEuzdX53bbvI4cUadUGBOqWvbnhzaCE8amdweIkQkFXnbvdCXi2
+TNFOzHHgcyVIC5Gu9ZgQfRWIJiv+U+/b38VDBH8wUDD00fpYGITcegyoo41tJjBxnBHbRWH3jx6
S0a+KVzJLO7A3X2ZRPj1ezewQlExWfmxwf317b1MQiIDFC0GJwoF5Ql1vwEVopLlVKOWdjT2RCFL
u05lVpZxCPfyKeJNZLWAoFrABirLQYeuLxgonkKLKgYg7uw9iqQ2bEFeXupYAjNIAwgyNGJ53USq
FM51JUBCSI1xHe1QWmr7KnCPzceiMzBb9txCsJYOVG/zKMDLjt7iwqTrP4BWz3FLo2TJoaUNX1Mm
7mHsp/xlUci5eXTdhfXPwwoWeTAzLmdHO1HuQu1DnR1UPWCZyroTgiywqBAopcGpKChE1Z4QFoHF
BnqOjKxB8y5rnW3zXBoqthrRSNnjyBWmdpO6OnbhAO+QxqKPJEAQXhKP8so1lC9qQgJQcgW0/r+O
tpemPsu8b5dkzdpFGvR4YSgxoOufS96X7UG2uk/WbMVOsyX30J90iAya1CndFATcsIELqTeAMS7F
/rN9G5mktXo//ClwrNja+26M/tE4FYU+GBdmNIdY7UdDVU4ocISeL1a0tqBBnNP2aHFuupVHUH11
5siZilQi7p0Mg8YPsd5MvUPtB8x+yhj75aDIo5qze5jKDmL5rQIxXSMpxosBqUkcS1ktwxn+3xFp
9709MBe074Tm00uGR0hgSnZtp0F6G59vLA8HEnnhyCulNgFmlnH6uvazzFEc1JehDaV3A3zJBomB
ySo3aySCZ6jyCLQK/c5RBF/PBq4H1qoqlgcr5rSAp9/9EDHr/0/TuwryFnpN6izqhyG7bgjYYW8b
nzCPiWJwy+05WSMKC90q/qWfDQ/von/xBnhRm8ZyCfMAdhcJD+XbRJulQVyUxBnQ4+ABwXtJsC+D
Q5jIuFSOrLElf3K4vpMgmcWqqPUhT2wSLvKgKyB2BYpHa3UjhnPzG5Flyn6iTwbAr7MtsIkFTTzv
b7vOn5oEQPwb729xfy/raTS5CRC/h230wnqTTpilE37PkJPxpSTg+Z2GHSDHy6aVJix6N0/80IIB
lLVfv/XtaOziO7M4/yGnVAg/JBT7PtSnZ7DfcBmuiLSFt2JouOlPxaB1ByEB1khbqgDwzDGQjSEu
kUyobKDv7xqls2c2l/ZCNOab3JH0PhysdQSarn/uG791rY3N0ZSdDgbC8SxhTo09xYt+kWjARxNg
yNKbVDcDEqi3HY5VuSPcIaf+INYBY1NMfJntMVGynPI6JldKv25KoflP+47AGUcJSgjNrQJ+A9SF
OIuj3ECw9zBdQBPvbXyhbOzIwM5J4C1i6aaN6TROUMBtQb0H0gvNeTAaBwBSo9eo+Efbm4eZjUC+
Zpjbz4O6y+gnZj/Oevl9HK5n4fNgS4CZWVXudsk/VtiJjQNTo3Ac+f3PQyvS//5qs6vXSfZNfIL4
+GVb77JPbyWSDBOlJ7mWCHjNuNIz7qfXLm7MCGan7v9WLeI5i/tcjde7K8mnCVNc+uCy8vKX/BmE
dn+9j2iX8reQ9MUHKWplSE51Ui3MbiXzBrVc9BmC+4ICZpLuZMP6baYHqqTEnx3L9IURJm8djz67
I8geISWcWcSaGbJk7DgyzjsoSfZOkKFpmLlDgdJdAhwRk2s+MfK+P2fCxpg6t3Xngp4gA4/8R5hR
eSHZfL5BEMyx8XKgtXpTSF8+1Oeeon+ELsf5Sj4ogQc20+iG/jlde2lbwk7M10x9zmdUOcWFXu/3
Q9U+UTaHAdO4moomRlF1eCKxMGoC6pBomZZA4gndeDVjWs5Ym9hSSxWdn/hk1ZOty5MR8h6GBygf
XEcsuh79ESXuqnWe8Oi2uc/Ecw9bWdslJqGDs5i1OkgOuaJkwe93B/LHBztjLbK5oCr78uTtvA1b
vYFuGm7530pYPmLccSH6nwjcJar6mcRJpOeBKKBTb+OMSaxOx0dZcfbMN5mb1JpurR7LNVZ1/TPi
sc3qOg0U0tkxhaEt3gh8S3QHPbns6RtOMZjk9XhEHOpCPWfBuhXCJesbEw0fFeEIn1TQfCOPTb6c
zvvqcBAH+wyu3C5xETQ958yWSlKYxeH9viBTR8XiHPyZMIsnc1oT1y9fzph9QkR5LxfoN+FEd2Eo
rhYK0tvS1rKqcFLzFs/dZh94azr5vjGGAVFA692kvCQI5dloweYRn9BzNWNlcM7XuascdT3q1U4E
DaEbNwfMfFCAafRBJ7jjweGK7jw+qe15punYaTr5bgSBBCgqembWX1T1IcE3D+5ZhSWWUxz/sJsB
D7XPoALadlSHTzHPMZXctUsZ+gFGNfjAQWs7NtUdrmq9A1QSrCGNM6cy7lAL66ji6rOR4A5v4wtJ
89qjUrua7QtQ9W6WCl2sTYXx5X7fT+HuyVD5qCmwl1ZWPIo+wJoo0tS6dQTr94j0wI2pS0SJ/JEx
dzW66AVzQcHjCumM8AbeZksGp9YS/gY9y1HRTytIx2JxSSLqLbjJfDYdyfTBtf+6SSVumE+pIxxC
L2skZ5ZiCIwvalJPjjimbXQUE1dOmIsHkTDGzILvD/Az7AeE8Yvubyy59JsvH2ZLPnmXIvDMheTy
xAUsXEqpMG/p2HVIqiLJfjD03ov+iqpfh/J/uY5pv00Nqus4gbSycw3/+z3epHJomy9aEk5xWrx7
tv8p8BpBiUFR298UTRGUdLBYm9zXibvn1OoqXCt02L19iFlmdDAebyUSUTURsPkX5LyUvRljXyUF
MDvq0X8+Kb7vWF7sWStajyMAp0tBF9P7O0zxUiT0vbmf/MI3Qu3dxiuII2zhNecg6UK4RIroH+Ec
s+WKYsQqqxJMASbtYAG8zVwnpyUjhBVxExH51n4K1efLvJLFw2weM03Dtaz1c1nt7XR016lh/AxC
LvfBAX2JMdPMB4FNclZu2WbIIkFhJXh4V10joaPWNb9G/R6wzCtdVrPr2XS4vY1JpSOfWo0stxNy
sUDhLwhIr6aEgPF6dvol7YtdAQADdv+/0PDGYz/CWzqUufC+fPudVfpI341okncl9Sy2+mxL09L6
ascwCPvYYj3p50+LvUtTSX4gB2UeDtm16EyCiudLc58GKCG5td+7yKCt45+7DVstabcsdrep+6Qh
ARYWGtdTdUsRc5D2JDt1NykMz634q0qFh1b8LbuEZ3hmDKPxNA6qCjw3ZTfLsHL1W7TdlnG+ABEW
Nnr2UB6uTOROiiSKkc627yV4YhEbogU4dtk/6FVQ1Gq5ebm0tBPnBOC8QU8o4rOsxJkhb8p6CmM6
SLwmBXitWwhpKVaPuT3Bs6D31pQTbCv71xtBPaVuKi1NmBmdksZAGog/DrrwFrs6VPobYTQXQFo5
XYB8u5XTOyXKWKpwYmNnLARbHzO8G5+nVCXm3L/JumzdIq8kvQ919lM849oLN9tFKRTqv0kY5oWH
oRJORY8tH1OGqZUuSbk8QJQdA9F7aIHeMPCRu+uloZpq0/sXjCuIh4WGJlfqJiKR9+OUCOZNeG31
ScjYnh4jOWUyJ71XOz7uv+YS7/Pm05xdofiP21c5Ga4VXz7w+oBZfSjOeqWCSf5e8n6VjZ1teKuj
ToWGiH9YkVIom7oERH1dCHEeo/rRUa8cshUggftIuJLHwQnWg1i6VxCahfNuaztu4On0IMf8Qsse
U61e8wdJRwVMAzWgwlpiFMkBBS+O9383Vhaf4AvUBIxMhiSFK7yUBuUjCqQA0DCBTU4CasfsXIxD
Qzfgy4UfGKQSEHFAMXrDao2jwdOyDUI6bfKWjO9EEpZhXTWxUEo2qcr+ZIWkbEDRMVf33oF6mrDD
xCEHzrpN/mQBHTVk0Z1lGBLJtL/0Aq7uWj3D/+DHAUXLMdrZbprO4OXZKZGYn/S2H7RVT2yE4Xp9
WU5DbFwo6x4YLSxCon314Z4pjnWTDJZ73GGfk/oaTHdqj/66BE2Gyj5omITHvRwHg1qPsIbFvwfX
Ow+AwqsME7DUcx8mzUaeWXwlW6/oiBchReeOpUXUTz7Rl2raKyb+e0YOq2iNrLwAOPIOkouW9kQB
nobfgJ2jNdaxWdDB8WIhexoFQksXLQ0XRCnAAg03S4mbsTljjqj3K0bPYNIOKjmAdQqTio3Ks/p0
EO3AbpAjGHzQNOm+6Q+4iTPBh71xRCVT/8g0I6llwD05W+YLS8Vbj9PS3cPgXEXSRyKArNFAlaKK
va00MKv15UpW40pzyw4RsujSuWdi2FWOzDoA+h/SLMsP1LlclBu8wfqgnFuMMhLkh/DaWh8QBM5Z
hWV1NnVHgxwSVRrWHntYyRxkZ7MlIzjESx4UCbm4lkc5+zT1wQmfzWYukSNj6ou8b83wdGbwpxCq
XpdOswVQ9oGcTWSb3lbug1O6sHYjtHTxhgPlGIt7M8+2FuoMu69JT4/cl+DndnqVeQ3dYdVzVYyH
u8CvVKQFc5NJnnw9OMxuzxjuWlVz5xUgmEkmhQF7oo+0uK2sWTnDqhxNnzwozYLQXIRtL227lDrN
ZC1Z8KIgM4+sRdYIg3pLIiff8xMekPxt3qFKpKmAU0dIN6ZEpQx96KHZBprU70SC7nae/w86bjkd
C0QnwtRLvTR5fWPNnfUGWXppX8jlxUERQZQM8VbJnJve40Z9Xp483632c7WIzbXa09oaW/F3I8F0
lx2GguQeiYjKYNQ+Xi0ORNrIgA9FVjgYSBoV+rFJz8M8WZxkXnzoEkxS9xlinfUzU6oF1/Lx6GkJ
edIjCLG/SzzkJffO+BfvS4hUUWqXIdx1b04c9DF7NTQguLd6XojC+WM/+yulSIqmLBvBu0Ea4KvP
Z8XnbcM+Fgz0RxCHbjHpcQBYibe5blNC3VJtFVknkxWDnkYiUQGvUdE5bkzoc1XHyfk5hNd6Vcpy
HCYBDVH5O56jel6VPyzk3gfsywkHEusEL1vxqpzSedYa6UU3baP5//zASwqj5xbqI1yzNmc48FRD
nyQckHYTfpsTdgSkcBeAVwrs9q1QhlLgG9Fk8wHu+LbZoA3Z4wsAtM0iXLjqtv5d5L9jE2smALE2
W/uvrStex9vBSxyz5V5kWgaYmI5SF097Wq7Px+1OUyzKai1vlNZTR/scrOlmnPpmcgdRGpdC5YVA
w92w2ZUK8OpRF+qrcVfjcxzrb+KuLReIJf097nWj+EmSzchiGsJezb4IYI+xJ1twgwRjLTDquzs8
xxkbU6JTh1BLQOkqMXXccM1vCCdbMiBfn3E5av5XQgJZ9snTA9phzBX3nFFjVb0zP7/kOnfYn8uO
Mu1zBie3UakHvYZYZt5HMhR1QnTnsZmf+Qd1v1lAMSDZKfiCVnkqU+suGhfJzEU9ym4WaOUyJiq9
9KkdKsxN5hV3Wkw7YpyG9nCGn12kRtOLLgftnnW3IB2NwiQaxP5Wq2Dgk7RvNe0W9j41gsb0fL1Y
VRHETkquZqZfzKr1A3vj6YeDgJ4PohNqXeRT7MwANx+YBuU/dWaTMhgQIHHDRoua3WdrJAg1C6Jo
z5pL4dqHjbB7PTOCUM39SY8tf7RAD7A52GH2mcfLAMzIThja7h9BTKpOAo/M78u2USi/On/ymolV
YBFajnip1cJ4/KOZxHFY8+QDfL9XE+QexSEox3yoo1hwE264U3EV/JkI3HhsYejb/XhLnvjxwulr
II0g59z2RPK5+1YRILVYBRzdNACSmhyjc9nbkuOEK6kGvephViQynYXLhf8Rm7P8UaMWBIvkh5mH
prVtyGtd7weDrXK9Bx14iU+rOOleyqPy+vw1FUKaqkHG3T68Hw6WjVKydrNFrfc1YbsjfYBDZOAq
eb67K9QX4FG9plowu7gKg39k3fTzK9C6TUFU1AIOtwK2C3yuWrPLnqf+AWXmTviLvYVqg5qkTOou
tqYzbyiTuHBWP2AL/80Pwvm6GPwBiHs3MDOwiGS0Qfp6fgf8Pjq1Vpg9FPx8MDcVD+UCLzxyN6+v
paQF0LNXqIA6gIoJlr8wSBZWNaaqZpxnXzq/UDEDUggiciRIciFcSlWc4ZlIQGfqQBSx+fVkTd3b
IJ9PoV8IU5D2aKt/JaAf0FrSfdZua3pAYQJ7v0pOxrXpDZw1/B3bH1AoxviMOoFWhPzZfAB62HKo
720weMKkyi8nrMmQ7WXDd5B6Qp26Njo9+ASW+leeIO9R4de8dgE75LBm/B/ZOO9k6wIrBbAaKF2E
WiGSs1drTQ9dBwx+QtRw9P746w/fcMsqfVNbLsj/B783Io9yuYSxKGucTsQZ1C/4plHu2qqRVavO
rb2oo35yHr/DYKVctxZKVSu9uokD+l//e6inBaNZ9Z9YDdD9o3UoU2QsVla1LAvgqrjIi4wyPZB1
CvlAGHJgsnC+oEBoM1itwjleLhljs4PEjl/SIBnXRaeNpeF+cwwDYrjqq4syK3h9BlyNa8WZpYcU
7IZGYooXfFCE8qYyR+/ePc17StOObD4T55cEVgY9pL9+rjfaLEUnl49SZrn4WWd+pcAbjR3eSkzT
blrcRehPwWsObzOFVlzhCmnm2DG/E88z2RLVY23oFdv7YFETDQE+luculrt5a11uzK3zvDwB5Ay+
Rs2tsoEcJZYu/sDFr3x9/ZxjUSXzyfkrvO2QdcD2A7Xe43xr2q0tntPNbXbIX15dDjj2NAWrbpTn
Y60lbMdvCr92Am+dlQmhGcMC0HzQd4vnJwi0LoSMKEFSEtWbNcnLTahFFQ242ucq1RvB51ad7zcn
EK3q0Th5joAZFHLzynUkMURUkkI3H8xKNeY2sVDGr3Nxu3bFQVTb5jxMMAsvJvUanP5xeAmyDshm
rj7vzyqkyR0MnPXZEAQRpDwjSZWGiSSNOUnVwGpitJW4UjKuTPb0B7o6Wqd1cd9UI33qeko2mdIf
wEIVoeDS6bddpYto+QtQvViZuVGhGx89/ix+LnmZB3FgvXuB8tOdIDB3xJaKyfC9EqKMrYfjMW90
Nf/WaSfm8D5hK1wV9Nb/jsdBjmMISnn3TEjlKZN3IP7ONUOorhJU7P7zHpndyE4khPSnKSieAGQD
bEKq1+RCsIJ/bT9ya5z6fZakcuPx8MmYR1GENS1Uh5POrKtITIfPUk4LANOOcoUU1126EHoF54Ly
eJaz8JSPpWv8DdvrL7nJ4h3G3N/nAiB407jsm7M5koy60RpmrqwYulJ7A48iFyT2dV67DB2y+3A9
0wn4S1pfXWGmeBFDR0Hnu7qJXEHaH3BZm9PeoxxgDmXwc9X166K32YA/6MLxhePyjNs88IOkv9P/
/VF/fi8QelcZkAa0jxWgdqBaYR7DJTtQ446jkt91k4a57UtdOFrvzP4lLB/OFGSc9fOmerxtste9
AK+iaZgeMg88QzqBQEXnV0JI1HuvQiWKurPyhM5EDEjyLPx5jgCFFoJWzWJbKhMojMWhFCAu2SJF
e9yvJo1gAF5Pn8GP73TH09j2TiFJC3m7uyuTeKRJuCuCOJbKrHhjRW9qNoNFbXi5ItZBQykYe78x
ec6TDJujoZRzVryLnCJYuo1qZA+FrH+xXOUyrM3pBUO8kY4Hc47SEjExBGdAmUuZlVKbNSSrXpuQ
pjYAYiguJ9YMdeKuTxcD0b2nXwl34/7YeLecMzCb8m20hZ+bACX1IVwqHVM9+t5uwbcAb9P/wurF
UaTf8Dnfu3MNserMOv8TSi8wsh2NpehIrHbNJs9dKQCvUuPOT+BkHroQyOt661nBeeymrM5+l0pl
5M+q2vCLwLvYqTxCrw60z/xMq7rWv4t/GriedEhTLa2DjbhuWnRnnWAfOGXao8Ve4HMYE0y7pphp
/FTc1KsoMOLm14UlnUR5BVkFz3uQu04oASpLwJo3a2SmYZ59f08o7oNW/vMqLuAC+P167zaRwC7W
2N3UBY+v0x8WySV/hNrNIVn2q6GVB3WjOIHE9t90IZm+Y9Z1U4gEzxeIv/AiTEO7dH/yvae0ru+p
7OjZ+tv7qZk6NatTZ1xsBi5ehAWUFI0zFK9qmM5I87tEHW9KswSaW+YP5stBMseG0kwGKv6iHSOE
FBDaFbw8nRr0+bJtzdz1449kAW+L2/nDBKWzGqt95+NQ4w+lYlPjjSJc47kFuZrZ3p/qmSQwSl6Y
BCxfb5C4y7Nk2WBBXOcqlkhWfVGb4v21The7oWh9UkCN9jDtfVcNeKgE72SMSfWOjuIbxSug9/lc
vBSTNS+j5nWFty4Ek/20JqaXV+hkDGvOn6+ngnyUBsTuBejBs2zDR2JR6x8jRbe17QNCHZ0dMSsT
IGqaXvPFGNE1UMh2MmwX+vEi53zhfcA46QlMu/RpJJVu8bmEG/MNGbq18kNJO3zCgrvP+7RKQsAg
aFiddB6OYDP8GKh7J18+FNqkoknLOuZ1ETrSxPSWFLC1baSV35XsBMbFWr2JixZ6mjkJAprIvDMn
0K1nTtTQMoOSCtRcoZPcezYAx/7oNAifs52xrqer1/gaNcNe+XIXo3dCR80w3lQ6Pru0w53t9orl
yu6N49nNAwyAK71ZCxTpOlvU+FJsd79AtuAhxxCYdEAFWyv/RsWKASo8jYKM3KNV4QCQZyKm9tlD
wSP4SPyk6DNTlYtmESFbfeTPoAPPxUcfjPpA9WIDwuSp18LFIJO6PZNhgt2xdPWWm0ZAmZB5T3Kd
IAbc2DWnFYXBIo5d/IoPxrUe4v2f2Li4t7LQFv8CJ7xTMDvAe7hoH6EKRmsJk5CFDTgo2QB0YIvZ
EbgLCZvLJsyHyXxAD3pBVcDD+ajKPAVN8qzDjvah646YZ+9IBcRaZXi5BUoc0/NmnEOxAqNk8yEb
6IHhZoRQbgjVxsGrtllYGbujCdwVmBV85fvvBGgtiNmsqYHenjpZWEfYniyZZTCYumaNtC2kMv8V
BMvRPrndTB0k88ax5Er7moLvM9jUSX9LRVkzL320y3Y7YEOzk/0i/IMdc5VJPRpe4H3uzre2Z3d5
hxLKLCWsmB9L7M1kf8+Ob5jNKJAuEsWIG4pqdB11xB+sNRGPH9EJP41XoG5k1wpSvgYkJx5VHXSE
L2uoauQduBizrHFi5zJVggUwnoiTx33CBRZhv1tX+g/CGQ+dJRlrU9Ly8Qt2m/hpXvX3+Ku1UjPu
xaJsT5pWnPo/kul5gMG9Vb3zD65S5rpXhTpiE5bh2WpZRDSEmwwM90xrlCGK1+hCyk2NIOmtDAll
eDrBVX9+WOCkE4WznsKIIX0TftEkZT+3c/c4KxZB0qWRnLE0zUHlJYo5IlNy/teosMvbY0fs6lps
U03caB82bgsbTqXRWbeZ2pS2mNRJ7blt0llA1i2jCjbMafOyBwRfanV5UED+yMkIsGbrGCyuRKvT
DXc0WVxtbJaw9Q34GTMiQXHHc6whsQ7QuaqwN9iPG02dm2BgknRAezIgEU4h+tJoIi5qifEeOS/2
ugjUe0OSH2f/k4LvVj/idp4JgfvKJUpLUpHCJVRNMbMiKc+NsYzTKetyLh73Ymjyfdx7W9rE+GEU
iOW26mm3g4syihgngMWag375FluiRRWGSIOfqab2QrbuuzutCI2Otfe0LgskoJL7YUyZqiUMsf5X
JmX17EtmOdH+zeEeGA5ll77Yx1hU/IfLZElsOX//DxcoAxnhwJ29V+9e7J9+OhoukOJ4sNYNlr2J
yl/SPJFg7ZWdxXYFMszo4OaVVka9f0Tnl7zSG19iNOFEa/k86rbCxxH8b0nzW6C+nUY71xKn1wuy
wEYxzE9yF/3jXuBRcS26bNiIPeSQ8i33sD/Nc7IYTBGSBly9d+D4z6wtZxZVNK0760XBh8LaN1My
NJjiwm4pLdF2Ia56wlUph4gbKY0k1vRQ/ypKJQRgVH22R8LmVGcePZFzTgVuQ2rV6GjTceeMPoq8
e2XH6eFXvYWNDvmAYV11RmziarCifOqf5Xr94IvlbyxeY1MzBLLbYCLjE8+djXn/oMud2oa6jjwR
WnvVlnK0ERGXxYxKOi5bdmqR09ZN2ennXqbkqToW1TSdvWdQZUlwUdY/9d8CGo3nftx3F6mfgC0k
ZHvo5yuPKi+gD1s0B9fJGeJ3BaKWkDdPzh2+asDNM9uacVMPi5mA+XCC6FlI0PBzIq7YPBXgzHAL
E9KBlaVFrlGNYxiDvLBUk5m3zvfo50un9jCcTdNkfxFQHFHMul5uCRY8gPJlDJK0qoj53k3aNXgi
Fq8Er0jSoa1M0aPnsp5y2lTXhpobt3u3ctQfubZB/Y5wb14HCrslSVHgBrly8I6mku2p2Ov0Aw6L
Xmz9TwtVX2JpiJU8s6OuWM0o4BEcWxJOSJeNpYJiKfaOBNLJTc7cbt1d3oKuzC+YsTNTDY3XXZ4c
q0XKFXFeCPUDPI+AZ3q+H7fB2SroYgB0mWlmHO18DMmHzHS2axTlsHwjAo4TzZiShGM5X9HmMzU1
FqZZS60vNGLWQyeuQ9jYP4JPmc5w7mkJCQcN2pahKLjAyG6XPm0Y4Ad1CucXhiNkUGl7N5g5SAJN
p72EhIhlyyt0+XYISuP+yNbcUaBbTYuMw2S1uL8AgowMGAGZ346cQN42I7lnqipsSfozVqgAJCAb
LVg3I3SRzg0nsWvN6H+cE7Rlq8chsg2l/1cijygojSiKF5qrKMA/JjWsBAqvfxej3X2u1fW+DPr+
YykiU5rmMet81lLy7BWteOTa0vmSXX4nUF8V+Es5MURTCrxXkthETuXz7QKcTRsEMMS0t1lCYUPP
091k7ylzzHpwd33Zwc7LzNMMVxqdDAP0kKF5SYauRJZbnSS374uaCnGbVDegPB+6Vat3q4NG8Qw0
RVrtomHkMaJQKBfZCOXmYOuY6Ztpnq6L5zD2YjNhSs4mfFF+F2AuNuJg4qGdqK+LzAyxLWSDYJyU
MvWjznw3KEzep696EpXIB8pmrvI4iausASgsVwAFcno3C/OBwssXhzZugjoPbNV/sF9JmQgXG5yY
mLuVYCgYmY9Prn2khgLKCIYmFc0091UR0ryDJznGDN57mWlsaJLUUKbkFIG5H9Mh0WASn7evQyUr
MiIpPEmxNGVBpg4QPBw9RkHXoKKIXFrog50V2quHyOZodCJpdqQVdWtdCvtC47Rx2GgSv7dXoATG
9WmWjCBrHO3u6QslZ6Svq/Z1ADtuBINt58+rUt1sjX7TDxrjNUcXq4Q7149gWBEdNm5Ak4Clp/QI
0NNhOWX5eCUF9oJPM9kfhAHh5F2UTaUne1smVpPlAIMSOdkIU8g/Xcztjt/KnSIlXntaBDz4TbHx
D/qO3p8ktCe0OYnq0KZvwKUpmasSNuLxavS9e7rfOs++Yb/cg20PvJ1F5RWsMCysdXg24bXfxtGk
VPhmIqnkMIVnHPbTRz95eaSpJ7P3PP9Zue6SMXzpgEuT5coq2hQ+zrNxZ4y0m3cQRScQEuOsLlN2
YlFZF7D9AcqYrW/zUlas+ARQlrvkFu7W7nWkmrsxErS5dgninrpMW7CTpC8dy9ttQbAiEKGD0m8D
BUjNiaSX7/2vm8DblrPhL54psjQOKWYODvsS8A6KtLgpCgMkt9P8+SkMKbUKV/dlJ4VbkU4SsqsM
rYQCh3CAa/mpzWMlOG5raUqdpQ+GvyAlMqzgweRa/+rY6gXeA5/BxSYdeuPzrQ83ppDi5DBOJaZR
IdaDZ8MJmPu+t9G1WxVszdTE8hkwD6wFMywI6SdyEBCr6oGuobew/uv5IiAIIye0ZnAYGq+9X7Dz
77bX3A9vZsmbJLvJzGk3fQhfuSGtAKOU0DjiSgdcWPV2l/e6lyl8G9GmqK4wXxpecYNROOOsx6TF
uoxLRsdVkH2ecyh4KWnuxFuxmWGgbXSOdTI4zO0FnQtmBWhI00tkEhYXU7bGBhRoxWHVpVWRRARy
ar799+ymNG8j8bknTSx3R0amtap6lEhcRu8WU0FcvITW3O34NqP6qshhrvTFJ5TVrz4QMkhTDIkV
LyaIvxcVjtTra6iaPp3SZZ2zj53o+9q3WoK/Wre7MfdvRIygtDwZDUrZ20/0m8WfwFuUyw1/P2IC
vkoHP6VuagxOZ8oVmH6pxXXZYipisR5bs46003U5ZpaQlfwpYGkrUA0y8F0bGy42nMh9ktQtCg/o
8Tm/jJx6IJZUCy97j1IasjQaSZVEI3gUPSwJspZRGn2Sd7B+YthA9X/bcCBWbipsF1KQzEvTl8D6
Ct80UcdG946yh7aceI++aFvgyDVyXLTsqzZxMZLfp+mbf+WpMt3Sdra6KEXqaKGPNDSHe9L+buc7
jtX+Ys1++mdIQ/uep321Z+b5p/2mFVq3bw4HqEQvF5PoEs1YaOvpD3Uuz41OaxBJC/LSJfVyVUFQ
197xLEtmqU8/YlmuZpb9kBJcO+sV1UX+UNU0CIwccWUtPOv2g1C+qi0to+HczyoraljoOztmSVhL
/4o3liN+egTR2erdvf1S90Ap7KmUO/wmepJtSeg0I4bGo8WW42flqH+eipGPimKNqyIVPaTElYFo
fyFVy3HObVYMQMT3t4dIsOpr4ZnSC2UOwveMILuZxDQEnpsE55sJLrNO+Kp0wSA8Q9UUv8oSKCM/
gXOk7a+uMKPeBw55TpKeS5gqfOQaEuNzeJQG/1M1pJ3JYM4B0g2A5CFIduirZ5EXm/7IKn16vfyi
0/0PpOj2Xgp+RDKBZmMk3d67RMunU7zTlWU0bgl51GYLpird+cVlahlIvmvxVVssRQWpT0KpMQja
hns+QbseY6FKpw5zmNaILp2VocS69UrtXiAoG2ZetF0n31VFoY8qQ8P580CSkRsADcM6GE+FysHO
OXvWupaFSBnrocJzht/HXAcRQWPzqbH8rUCQtuOBZ93U50o9tWfIIG9FZcIKmIoHlwglECfK5up0
Ee6ExYFD50y9dgrzNeT/46K3rGiIBJcIGLhG4dxApfh3Y9P0JwNXJxV03XhWhLi7rS1TwzhAi+5m
DsWAL9rvChr6GRXjZ1eV9i+auqidivdkpVr2Ohv22tRw5p4onfPhQK7MzXdOMWpbiJS9C3xsJAzN
YIBgLM6e/t/ZvZJua4fSihMLmULv7kDrYgU05x9PedTwjphQyNr4GJbCUeTK1E0NWV16Jrl8qEJU
bndfJturKzMVmtsBMjipqW4vYm+womaMvW7XhC9BMw0TY3USWwhfDqw2KsHaJy7rToLv8Gp9idlV
H+NGGjx2ySurv2bHBAp10ABjrW0RnjZtqptv0F4yUDFU+cvGcNueYg05ue1W8Flzp2iFQsN5egRy
FJsawpDgFTgwxXLW5vDciLb+tHKXm/Q5Asx421hBO1iYfu8knnjRdvaVDRHT9JPhXGJZGZ2iMHPV
DW+C47XYaWRZ9Az/bhYzugxG4KQrfMUG9QaPIQIC4piK284KvgCFma4iBJtNa5R0n4AicesvIlQz
4gm3m2Zv86EbOeKXoEKMO8wRzbQ6whCLMbCZ+npqu26R+gkTE1Rslv8ECcHDeevCntBb1hsFJ8ME
mWUFWVDu2GpelpQ/+ei4gIIv2Ec6F8QPItivPgi9ivmDL7OXLzLnf24R5Ym3/HJzhS+8GKWUnqCF
nsXqIcAu1nf0diM4eX0wLCvi911OmpWVJAQ9NPZCqmvbfoPX/9p6FIhD6I4jWEUjGNPSQ8bA0hCZ
AZJfyh9EPSfi4VuqX/8DVPD+a/xFleL0gdtOCTloaR5/3U+ZIprMC8R9Xu7/SoDcsBQ4H1xFoYRo
Pj9jn6JrVyv+OqsPkgSwbvtaO3e5iCQtXxgaGr4U1PkeatwiUwNx9BAQSoSGVEkaTVPvjBldes/E
uNmkvyqI2WL0qoxunyQ+90bVu8pbGYxDMSivFAfcnWg5aiOQtevQcQFDO+kJ7V5PQKYHVasoweNL
+eW+Zq58iPcwpCMphzFL8YgeWiI9uQuqhHSU+SmbgZ5mDNRNJ2ps29ZA3a2R8M4YiVdPq0ucPe6J
gT9ZVVu0RzBj8vB7El4+QmnzpxIX43lsFvrPYm0tHb2GmKOfGNHY63GJjC1xyuTEgKopeErmOlx0
YLMLneRASCGl6QWRgzcCjO9+AeglS2OPSLlBUe6FAJEMPTPAfGxELWnUjEaqSJuCOk6nVGXR3bJp
I9DAe0iTae1NQDwz184nhEQRlqPD+1Zvv2W1gAJ9ct13vbUnEXI5q49bZx5GWBxuxsLnRnhkHxD9
Mm7WKQbyhwv0kKjL0/uwiXmmsNhDG+U2fO59ceVHAmLExrqgCOtS0QTRe12LaFG8j3NFn3FBmBex
SN0/QXCU7FY1zgmaGA7ebp/2vtaOTJYevx1eTJ4z6ZuTFIa74G1lhw0dPinO0RS2k1tOCzGGd9jM
tgBuNr7KpCED5njoGhdRpGn6dVc7lJKVCMmMgg/HqPwYryVgahmgNcX5VaxNOT1cU6aTs3mASHEg
Zvl7cs6RWPNkfHQ7TChPqVWm9NHPhQNebCmzFVRa5p+f3wFZfezltEhhmJzaYVPAMsBrKTjjyuHJ
mzd8jgtvbDfu8aCxHjdSmvQfwcbLHCnJj8R/ugcf/nLTxiKF9d7/nFSz+69NXm6iJ159WV2Xdyct
SfdLsTidCc81p0Ygw6zaKlOuOv8qtbs+3EalorEXcDWeCB5ZmShAc7MuoL5YH73nOBn8y/wrvr+B
EIPq4+XSB7Bv3NpDd779uH3mPmQgdqbfvRCzwtDsbkMC97QW1cteAryl/RpXfxEDReArZjr5NaVV
qZvaOGbYQQiXQucqaHPAygjs5de4aj5PKuJkw/vebYBsjMspIDe0FDEQSIdlWTkZ9+T4qbw8pSPy
MGgT8+QRke3Pzgp5tbT9k1Js2pmy9FyWOBj6BL7hjSZixbr+qLlptWOXUws4eiH7s8dfxg2U/tgn
1k+7WaK6eCn32MoSJCMbhZKxxMQJdraJmMuiPVp9RMO+dE2QzYrBH6BaqXGUpPVON5Pyzi0VeF8/
vgp+qlKR4ybOPylTZYWE0huNSI51vuJKK0hJ/kL6mi/9Jd+4zq2H3BcmdJ7SyE9ly9EwSdafRUYl
62E/rUMlTnjXGYuQ5oef7BgblSu2G3TVoGEgZqolX7QZTdYmeQw37M7P3Bb3WyqSDddqKlbC+dXM
s6cCEzR2UL1FHA+zGMVv9Eo5dGkvoOtToxxIA6S3mRo9jQFNXisDxgwEwWA9rPJ/swbNODvhgWEU
0RvE5Blo/49WI0r0gSuOUuLl+5obDwVkwdG7PvphlRPxyEvLZU7h4MlnE3TrE6o9VUPtEcW16OsT
FwhuoC+9zV7M50gM9b/AxSefBH7bmHh18KAlztNIgXz7wpol3LSXGTeMjxxgFBZnH/WpCFd4TA8l
yCRU6VwX1giD5W6xzfxWfZRwa5Zc5m7d2aWYjPdVy1qwaT0aZ4AlCYViIwFLypHtSpV03bJ5z72o
Kl5Nlf1bw9Q1kIf/eN8WSY5W7nMJzfzKyQo8DHMC5lFt/PkWSNQz2JKoxPK31GKfc8PTAYu/0b7f
FEhNJvpOoHDiP90ZL3be+IeVw6JObye7xFA93lguYcdwv0WGc+3WsLOX5A2LXUSygle0HRhAhmPE
GM16eSmSXPmZuw/N3A+tb2muvZDcttvro8V/Ozh/PqNPrtirCtnooAl4fwi7g4t7sGx0wkZVe0i1
k/hrOSCBi3z4Q5HjVnOKYYbNFuKTSJOEQyNoeBKk4cC/UhO5Ca9wpdk3TQqCILhN3XMFKUY26X62
NOpIZFeAboIpex1TlFT13oVkqJbIPa8zelcXNSOXTPxn2qFO/ZFnh991t6Cn7LleQdSbLFbN1cFK
wok2ejgnWMVSY1F1T8Tbupmlh79oOXMvAwnaAtXS8boATEFLWEAa+UR3aBN932RuXkPb0lWIDmk9
KPLL/YiwzE9wmWcXiRRj0hN0cgYEty5gD4OpBydxNWGt8vodAzFXVW4gVLlGOyQQ3PfvVu4JjowY
u/3FhgJNfspCbiEUq2OM3FDn0n7sbbWFK4HMTRG3pnfisKguWJ+/scWqdJpb6pTlvVSOP/L7I56A
u0Ca+zCB8rvQvBPFyXou7MJit25qBgcAGoOmjLLdKz5oqVMMEz7TwGzt2rQSozbczN90wwGbmacu
5aZb1sk8NIAthHYiLVgtyI6mRvoWupErGbL6kev0P+v1UtPK/W5JRY8ZGmaXROxLqEOxMfcmQB4v
0kBBEj0C3fqKOu9DeOGlUzW3RhPHUJcCHdPeCZFraBMc/2gDpxiJcdRuQhFal9nSeziIdO+p1GKu
UM2VrPnMg40qARGMgBIseHQyVYfnlowC8cJHUr2dD96ex/p7gyT/Qx8u/xRbtFsoncyG5RR1QDyX
8c+D1YhZIvXlvt1f+0yDxmWSyGc2v9bBN59j9uKmNRcClwacMj6tsHSMQ6oNLHV9mNooliefmDMy
MQywxGDOdWJCP3CoIUA983fCrNZsDBW53pO3d01Iki0vgeeAxaygZNg+7ZVl1ByvBaW6NWIOM8Ff
UymONbxzu0xkk1CVOureJ/Wt+J15o7wujRzt8otTo7EP0QyMw4ZgzSRPbJyTbIzphZUrUNwcYG/d
nXCu8fuFVSL6zfZcexrJf0wZf0b/pm9RuFg8LM9bm2NqdNC/EYUCczaZpX0CldEUGhPiPBPIQRwL
muQMF17HIy4kzCMwAUP2j9aGXB+qIZqiK9K9NCa4Wj7EwvSGzt5pQls4qcN/Cp16h+Fiq9ISI2jY
nJsQmpxZKGnFOA1wMAT5s4pdpn0l6b0vff17ZC9x0GWB0QwqSl9Pt5tMbZnjtjQCMKXY5wP+9kxc
VUxkgRNuASm8mItcTWSOdwY3Y9VEHHH3hcelY49jftwjYURiK3ATedX9DwOgTaIY1yDFolftjbWy
X5ecOfjlWhfOA2gFDxJPD8wFPmCtsylybQ3A3njJQp6nQb6bZOj+qxe7KZnrQwrlO0hQu60vKHkn
xsQujbaCC42CZ2K4WxMTf7QARTvAExMINnX1Jem3mwEJ4xM9W7+Xb9cgAeZXA/t9a17cyua3yQzg
/l4cy52WxEKimZ/1WRC9SOAU9HUBAoBsScE160Bv2rqxLq2pOAlSh/z+qvnsB6YGYjaOVt+UevHY
VBAM9hWNzQqH0Rpa1NlkJpNdkRAa5fju6HwhXPJwcBt8HCLhtHq0/1bVjcl64MDgAbaMMonwVPmS
qxal17Wcaqs+VIEUIsj+cIRUl7XqZNSdPkJtdwEv+SmA6PmkemE0b/JLJYZ2EqZnMu6ytvYNnJHm
qxwuUD1zpi+R3y7blQDKzsTr8clI6qLUTdRMTSmTUzSbniF9j7pO73k97jiaJJUUknTC+/p/YLN0
+J4WI8GQzTfNvsveS8xLhN6Blcp+V/dUd1szMxEv2vZ9O+NsNu80VcjUnjIF3/a1eLwZRC1KveR2
UmmLMnCqoz2O6aBJS+WCTaIsZKhOThp2561c6rFACJkQVqoXZU6Iu5jqRcmn8SJ23c9HObKwDjws
0CEHW7/wmsQiCBsQQ6RuQihMiXkfazUNrYlz5sqGaEgJaFVJgaaYkAu3aTPfv1/rQzJdpy8DGo2F
rtt5ckyJVDfIMfaE7Ec7x+S9+MhzMK4oXQsUtXBlK4wTLxXVyac5tuOBenO7+lK/OMIOH1ieBuWE
6tCgaUx9P8wJKHwyMjpr7Eq1nxeY7+H9FLMsnilTi2FYUG+1w1hnAx0/q2fVX8UnBDBawtlT6zpf
p6UFtpi2/AvmhjHJc8tvui0C2lFTL+C5955e0dXsKp30bai1HsHQYbBXSTaz4NqBO9g5gmaVkEib
zXq4+WpWg1pUZFALhAjh2Eo+4fuhcw+lJj5HZHcUwoBRFfdu7tVEvbVJDoKzXzmEwNDFQqFk2Y4O
tVuSc4jM463CH2zCom9OK6z36DZT0ZfHMzvLyznkbKnKTfQatP9QFa/Le7cbHdICAj7CeDud5T+r
LUOzcLz+59xQ1RdnqxuEXFTZdzpfPengJt7wECsgILlVyT8r7PGIsTzSyD5mYhgpAHcRaMa8SUQM
ZD5HeovUlSD9RJgisgE0zZkIdJHraIZREkdlUYABrQPvWduvVXrCHBxrIB1Z2v2cFonUxfb5P8WE
1V6fOoMkTvC55F+mWi9nEiQMePMP3q+T/7EvL4tFecSCR4RWdJM4MS/MU/2XBnioV3X3eAHLWd0q
QcGcz3MrPVwgoSaQh2pxhDZxFHTyVS2xEqpdSDIM8Yc8jVJZ42GnTIWz0bV6NlEqVkZCZw2YrvpF
BxdOG4+sXS3RSKKu2waN/TVhx7LEhPhPnSa9R2rMmTDRtStjCE4HoYXopd1U4/o5ow5fX+PaYOMl
qmBs28EVg98ewqr6Gwk8e3W3RpGzsFU9GscvM/u1rUQs2Hacl5e9vjSaijjI/qCxBnEwrVlpuAna
DNIms4Mw/dwvQE2W30y/OyGhccwwxcxbQO8dhU7EK9PeADtW9mTad8A98pC4TqfjCXstwHqUQQ0W
oPIDkniBai+eEyNKW5uQyiJB74Njf9JUvbA0yB6chtekP6CuupWNqvZvHmblycXoJbN/tJQyzq0t
IK4DJMtFGA7Drirv4cq8xSHiYInNkurorc/5uHBVk/2/t7YwENE9dBdiy3yMiXN/WbSOLVWDniMn
a24Bu1PXTVhNzVfWmBO3WCIexeWYyMg93KzbxL4Sx2S9LC3PBtIHaN2TDJDphRafkJEKC1WnXR2v
ehz2ASKWc2OyJL/gRPEAPK7y6kDF6M/WZTGlfbY20qPRogALKIAWHmH3qzjdk/N9LXN55/Nqrkcw
KWkIoaB0M29IBIAygkl5M9DljDHehA4N0FOEyXxFmtwfNrCSYs0402BYR7wRsfyNyiFMbNl3rrDW
gDOxLI00CjExV9jf/yPpxD+UVcD17BOgQKWXGfB6zFd1WZohWss5Jm9T8UUjgltzBcArb0EkhopV
GG5Gx/RUtX+kOFtPTNsYKnhUaI2tgLqxu1td/mFpmE0RtjzSGZfR3x50+uqTztxjCdYeF1aTJKsB
yGmSA4xuMaw02TvNOncY6TAaK827iAxHBQyHX2wpJX6/72Kv6d278M32qGRwYKso52Z4MSHvkpKb
iM1+KXXCDHdd+SvXSuTWeHZH9nwISmKzM0kxUZf7ut3TyZmLU2uKiDaA5h+plhAJBRYTCFeKzKx2
szKjEpwrVnuggnYEb0CfFGBTd7/dwXMfnZbT6ycZVD5aJEXE9Wmjl2s6yi3PjWp1x1E0MeKCtoxc
cbuye1EO2bZrR9opJ4S4Xzg133ECN2PISSBaXFpgZTZ9+2nSmx/hW8bpNij8Wr7ISSz6vvjucWFr
XiLPsZUYiHkYjSTYLWoU6B+urZiN0VGxYQ17TC04qqzEFxu3JUTrM4MO7nqIMmom9KFvZYVtFnld
mNPslLwFuBXlKKFlF2qPnNk0CNG1YmqxSLVJw+4FIiPFKAv0LIF/HGC/XTusW7ChXOKIFn1BZHyQ
oGiuU40dso8+dPCu14JKkfiV2fti5KR2T9Tp2OisL5s63qxDFQdxF8WTwafPoQ9h1UKLWcNaPdNd
vvO3RT537Zsr5Mxh+YG15hIVPuYdQNGaXXsGqhLUnmXsjflGW20rWz0vRuI4IS32PQOpefPHnkYZ
+1EYcHlFy7YnLrUVVFHDYjA0JXCWwkNDiqkNpP1DiW6Lxk1H8wkPx9SiunVBxlUreE0TpREath+N
VKhSPrlC0KvIZ8kZorwMpvfPsPEu/YCbbIu5T06oH1667e8asApgPbsDmeoN0sVixrp4z+XOrk8E
CEQfcGaMDU0vYcExqe9lJeNfkVZgt8pKGsDMVQ2DL+v+X+SmcTgmJoAEK4eY1w15teu8YHzEVvdY
78Nsq+11PhwlWpH2byw73rtTVVdbbTp0+EK/8pMHcHo2JWPkqnlRm2Hjc7gaJ+qAOQInGY6/qVwI
BTIoW6Iapx2BBIAhxyuL8tGoQOePtuHHPIY/Y1cgSHzH8fnCBM60lBsgA7dxeV/PeuoIA+wB6cih
tVY8h8YmodDpiBw1PYbBECyUh5aNnUV5mcLoZPM9xfS4ooaKyb1ZQwjr8GnC4sV+MeYbuk2MzjVa
ZMRGcEZgo/f9VKR9XlZR6FPcBpipS/Lw0jXXqVv0lDTGhWUEOIfrDBFA9xe/3RODU6YmsJSlnYee
NlhUEfY2VXtkg0RS3ON42YRliEFYtO71K3GBYwWtT1N1bC467m+8BPqGUWimbkDcasb/VyOQFfg/
g6LKGKlSvgb8MG1Vr0aYTDk0qYGme5MOfdeBW6TUeI7+g9ZJMFvXdjI04kY8swJMh2sfVT29eXJS
JJHtihCxqwfg3xg37qJuE4JuUlC03ZQ/Xd6TC88Lkz1XO+PVz3c8YCLS0I8KosYnwoMInCXlYA8X
rvT2maLFAy5gFq+ylKKYhhldrllhUJkyDDYkALC9LeQl9HiBf4+LKZv6x1GNYHdEOBcMv9mpPJ/1
nueqXEqJXmCX2oTrA6IWQerZPGGXyv4YULz+RNYY1Hd+DlsJFCJttC9xatY+ij9Y8W6StwW8lFw7
oQfNEN0puJDIqZrcKfJAfj/NK9CkSiR+ZYg2nx/Vzvep5vntTrNtSmdpA2idC8FS7ATpQ9xqgvxH
P5auAVDGaZTk8C3oOT1BP86cbMLCPj7Hf1dt9CRRHSZvqo4/pMZWYIhgMc0kzrYbJNWa41jIXA+s
sHI9twHUrsKt/lKkGsIDI5truAb7s+8MloUwDqTVNGET8k0oFsl56O5+kAJiNEfiBRY/kzO5Oq7I
QIOo+9rRtrEIQNIBDdqnDRr9Dni19sDvCDbLf0X1dzdyXf1sRLqp3FKPuyX1lG9DtDoNeyacjJWV
YxLQcrIX96rkov2xZObZ7GD1s0rkIkHkwSNB/SHZ1woVR2dR7kCrCkxb9FTvL7RD1ujbrarTG0OF
YPC5jCTKDeHwJYz1l0WSjnVPPLTI0wtqH9AD2Cfxgi8wBisPuqGDgQbpaN7tVn7eWqRwihtJcM9L
D2XC93IOAbrU9oGZROGD5b0P9E0jf2fbfaFlfR6Uewse+ynLscoxULC0VhzR0WlYkY4Xnwcr51BJ
AIE0CbQr3klwepegiFmye7IAcQFARlCW8t4tnCfWqdmOscN59XhqerfvHDA0fTRWuXFjROTYTm/q
fg7zr66Rk0o0xODOTr3OF1BIGS8FjHf3VO3zly3w7CUoGVjErhAccsultDnvibFmbmhYtMheuwnb
k4KErhQUZ3A3zAyj+eODcuTojgxVTryjXxTWFohzlGOVy4jPQ3G9Z8UotRNhTDqm9D8aKGIWQLg2
7LeEkA/Gr5+sFLbLJCCzHDv8NHi2sslT2UIIvrHPZz2rhpTGxUXvQwsKiasLx08qAFfgdoM/Kjnp
RLd2XUd8wsFEMwuLCkQ/eHNAO0rnIpIw9GzQdMhYghErm6Sa/ajfS9ehwJUfZPGdLBFLxL8ERhim
rCDJd6rm4mVqSDRJlt6xf72IupydpWnhAK/DMFd/l8DEnXY0ENJXUNeMrqbZ2yT+za/npFyQPcB7
F8e0EaWvMlLCzJEVMH/x7jr/W/8vjjvkr7uJaa5L7Smm5La1LhCfYZxv6XkegXjw6tbCjlH0ClgE
AKhkMdSmHtosotSQgALgfUJ6zl0q3fx1HT0N6fwuiInqait+f8MsTk3wOsevghU1+IszpQogTMRO
cI+8FuGd3L3K1TuGiKxk2HrlPg/tgZodjzPObIvIvEfk8mZs3Uml9GGvX1ErNtjugZnKZQMD2e3+
kyAtqjR0YjkFCwWtSd4Y5uCcrZgvC/nXPj25eSoEoBH7Ujfba6DiH2B7rHLk56S/30EO2VUyCag9
sqJC/Jk5kxaeK2Pa5s0bSbnZeIvDUR/JGs0bbxmfMOiRgy/SMbl9qHmsiXdHNQ9aev9i0dgSTg3o
WjXVSAbGr10xJ5jsP1v/IWYc2xeA3ZCuXXZutvpwZ9vfzgO66rOC32LZiOM8BEPWYU9ysmijh0pw
xglR1jTZeVwNzfsVLvUfiPnC5nP9Wy5zdBr8hIxrUJ6fEOPA5T39VvlLPo7//yvy1Nxm7GcqP7mE
/gIGsphJiTGxboK5iaJwb2mE4b1/eGxg8UhWElpDaRuCOyDHSxm8CgH43Ok19Fx1rkD7/orQp5rl
yoGXgjrBAqLaQnHi7wV5DVTdIUpdFrB0tq1gDo/HPwPf5MzuP3gzg8QRvoV9FH63PLVXwrvkcunu
zwlWrHJQsNxanTYlKfNMIK+xHyuql9WSR2adoxM+NmCCWPF66m2BA+UO2hx2tGj/rQGXVBSMpbKG
70hrMoa8Dr35ppif/pd0T/u7BreRNSxEmGBo9qurxTV4dVf1U+eft2AJLAgiV+6F87vczdiWsY8I
kZY2XkqOsKe6kPKZo8ZVHxakO1Xq5M+zWWzWKd9CNmKXcJsuXAlrWLSpgGrFCw+B3/SuqZW82udT
ygG1CTDOSmm1aKd3DfoaAYD4eDsUXRjHJu83e2LTA0WWFMIih7GOLguPNLNPR/3rzCYoYEwu6Zbl
UtfIRfBL3nLqctCKKpJ4gg/jhMu1Wb5Wea1mPO+kqZO5BZCxz9raDuKptuRejGvIQta7htyGeR4A
cKmpiEK9pqXSiAE18PYMSpLPvX8EQYUJGXRxp0+vB/t4TapeybfW9a2a9oQ23dLYQOR13coeg31a
U5YMkOx8d796GGaEtJwLVJ/C9l8rGysfO6N8QjwuYu8gy4RFkZPN/ZiDIlRlf7+W4NO/352f68Qo
NB1VTdMtiZU4+26jWeGi5wwL027fHNiqxtouuzsKJZc1/pl3a7OIaaBYWupAb8hIlUc5/686Pezk
ejW+c9kpF1Ji4HJH3/oCfpkbXJbYperCwm2WYW7axq/3lRMhzBzakUoVLP42Od3NzTFPHQfSz3tU
N5blaEwmJ6vEjFH/nKXMb/UZ4pR7g6HXbvrKK1Wi0iiATf6fCYyS2x7GCI1J2XasBnY1NY6D2YOI
zA2K9gvXn1SBlEBiY7k66SFehHSDwAzSoDPaG2GkGIRSyZzTUo9xACwocjU7HWMLCUK8GTzyexda
Z/QOmvAfmkjt4mGx7U/iKrY2FTQump3+ZrRwjWufDeh1MkbeLdeXQhe+CgxDkYwFTxd/cK3MBN9r
SGTvciokjS+DLhCCRzSMkotKQEQ+6PcIynefsn8rkd+Sxv7x4OzYIfcqKOVDhlsZC2Zy0HTlx+Wd
AhznQ+L2fFfJ8rV8BTdsMqIK+5CoumO3O16vXcjd3TlrTqFs0VdMzCH8lR+0izdynuM0Ksf6kb9u
7kg/ZLSLICpPgoIsZuc2NicYlJK8z3LK+9y0SqA6WZ0uJ0HDK/XgVnbJoTITxf+Ti57gWKyqzHg2
SAnMNHUl+at/2TIq9N9JhzVa3AWqQPOPinJ9KUX+jisHGUGtGeJJxg/nFfPZjkBbO+vLdz8RzLjU
Ppr3wOQhP39JxzCQTRL9uoL34e5SZSlnJ08OGbU45OTBuHP470kDwKnWlDPe8jY3wyNw0G0ao1gk
c+leT4MM3ctjeDDtj+c84UYx9moQOo492XbRP1VcYaJdQN/TOeGx1tEU0I0zjBGTyQHjXYhK1t7i
qW5b+j1ELJooddQwgMaMVqHbBBUcs0UALcAFoHGniNPKvs2ugINHQHk3JIxxmj3vepC71OJ8Jwl7
Xa62JbC2drgklPn0ei2oJ46isEpglrjINIj1nBJpOysXgumNxDYBEqb0wqHLYsEWrNI7I/z659G2
gEApDurWI55YyhEfh/tViZTAwh2/0y6WwsYLnhCeeY9KwnVzPtq1LiNRIuhL2AKcdq2oa1skfDK+
SPr2dGntB4ojG7sRURU2w+ECsgFm+ApsD/JI5zzGgFp9YY4A7Kh10KxnKwyyKaT167oh6b4lp9E7
8B9u7u5KZDh1ogWDTK04+VS+qGcLMqI1xQ1r772ig3Qt165FvVrJPMAy8Io9atK9fAW0BK51CHJ6
AMssWcR6ejqb7l1QiATcMUhP/2RBgg4H0/se43Xt4PDce57Zt/c00dfeo3mOJTvgrWIG8NyNLQ5Z
ARjXmPvV1h2+fM4H5K9bAr6AFqZDF7i7dXF4F6NhSzHXWrr5/W9jSJZ2e3HiSmS0+6WrYjmpHSab
Iq+9PZWkSQHZevozmXW8gIqaqMngXs9hnHkRThf74/nJR5stikI9CSVI2w0+sgOGeTcV1RL5XDFm
hLjPMAdEyg/4oYJfmSDACBtGF0c7xiO2W2HyZHYLM8KD4pmKYZzzzsh9N/2SiX9wtuNpsZPsl2b+
ygu4ps1saxDUVKK9LJDVqEnsFDFhqfgMXhirPZDsy1HwPUu7H6ziXnowjXOEcB45mdYYsPS2kc9I
WVZMYkutuKYW4fyKNfFz0WBL7RuHpZ8YYRgldXXAcBmujxHPZ51qFbQkqnUBu+PbfuiEQhrDR8sP
929YKLPrzLTpVRp8b/+2rj2R02Hr8wJ3Ekmq9UuxDYfP1CqY/kQI5bAokiIsE/sLZ4aPPmqsdWV7
LlW/jYhXXrFxOGrHhHBCZwSebz14FI79K6ywz08RMtuea+P9h625aldmtUwmp7bvsEO1JYjluyCw
WOAfy66W+LF7hwMvJC2FJLQAny1LUzI7vfEbwRBh/1V2cohmD0OjdQZlKFAsIBqXUfXUaeQZgj2R
8fjKR4GOKvcZNGImJe4pomPfkLlXe8fT3yXzhhh2pq2MkytSDkQM9tDDA6xL4428Agtq4jDSLGxT
TS2xZ7JmTDUtz/xSfpjpB7WA0lboGOjZYb8LReyNkEksYyxYZTwk+OkSNn5FEqfjZLL0+3jMcJ+h
qcER2+HgfIDYE/FZXcv916cfjZeyWhrh/BdFK0z+NHHi3jRzy7H9JW9rKwPWD2fTffJhKBoYSn1L
iYwvOfv/vbxlsRzCI4BBgQ6MA232Gf6cn3IWFm6qGaOF3vAOePb/3wXeqCU1+XGDdBRUf9GpJUAZ
KOE+hA3oDQNNBWoo2z1ZEznwwWxQa9wAgj9Il8s1BjYjprNhxi91c2Vts8h1XoeseaFpOtGyO3+R
aHD9zeOt31Rz4RWE3nvhCZ8+2T9R7+BMOvy/OFe7MqH1MMrf1yRJVCSfapuSon5flZ/cJp3jsO8P
TvSs6ILu1r7VAHEG0MOK+deeZfNNdETD5KAwSxqkbu4AOSsV3HyyK4oj7ROfRB1HGpOT8uaH2xFT
/MBh0cMQTVrGkE4sX8iNCxb6PvCXRUIxBrl3hn/yST5copYDODF2Lr/pEPIaXn9W1AvcKbgtK+2p
x0Ys/OXTdxD5CMRvj9GAZjY+XxxXlRLTsz3ij6lRC3jInkZDV4YOv++FMBAzNM4cjEMA6TcJh0/U
Re+nFaa1LGmfD6pYhsJOYAXug0PCmT7vYVjZuNNUW1HDR7iT4flzVMZlXXpm5h/MmFcehGqFkIJT
Qcvoyy6jhHLHapM5PcJ7snWrsSJ9yup58eSH0Fdc8JapiEvOvqJ+eDhywLv2v/JERy0/tS3EhO6D
z7wt+awJoNEWDZRT50aGDrXTWcAsUAPjtJPJpkhI2GgTjN+p95jB0bG8ZQzZHdAylptD5WVzM9Nt
HXvaA//kfj/u7/MFQj+Fg4XvYlLcX2oWJaoPe0hyWciJ+d6Gl/hVR2rZWuuMmiyIKeTEqi/ZjUou
e3HaGLW9gr+qfHbSakyJ3d+6TTcQYaZPN2kiVhA+XY2yyYhBFIt14DQITm5w7e6L5/vXVKe52vzN
eVjmWydh7wr4UFbZplS4uW2DXSHVEzqHNSNIHxl11KxODUAgi5UtT5VIWdhvEhOpCQcr275JW9u9
5hggjyrX7DMgcO4+rjdkpD0Cw3lotUADqVDbCtfZ2JtA6lrvw2BPf42/cZg23hDFqcMtubolntkI
8D8fmN3CDOevoE94cYjTvnFBZftpn5mDQgSIdEFWTMJ15qu7HeYzjMhpAwiwXgLDg7CJYnWdndED
dHCkWmnKfPh8TFbghBfWULjRuCHFrnzanD3YbmmxZDkkahmJ6YPVyJLc6cCGfoYBqCqZPDDUFZ0l
ulUdtWsjuA9uyYVXm1tlgkYDUB8kqDtZNlbFZ99+ZLM5K+BGsCZGlHC1QJbUrFwR7yKleMJWJ8H7
ZFhx8uNwrxj/ZsOA2wMTFcVs++Gc7SPtQkI4yM295hUKf2zGoXvkvG2Hwn5qL21ulrE5BfsHlcPA
0VlcfLKrD6zHHfRZ3AjmXFrnXxXcykUXneuToBt4qPqS/b68m0Ve3qCERp1tIr9erlDcgMiVO2wo
VlOSsHYaPOGUtnNo1ONW9AGUuWKoZXnBDOUv0q5uRYAOU585MgUb9O/ol0UM9T6D+kjF5YJEG+eo
kG7beMQi0nj4Aogh7jS/0+7rZ8Z7lyUMKOnYhqZr4cnBqiNZFAuf/BIR/odH5WfkukYOUkL2XgGs
SK2h6mWFMvpxJDcvwIkIi7Qk3fyfwd0Ycj4ly4JASvXQKLxvb/oxsqESQ8a2KBk0M0Zmm+kCH+XD
RAVtbFub0CgtDEw0qrqX7fbkS/zgWIoUX+ZcH4OosHk4jtEAKMbOiY0o1J/byud9goU+xcLZmDte
QM6+CWxkb5feuNBWRY3SrkuhdNUFwbUxO3C4n0p+DU+CFWZ6HAIhuVYmkiHGRmiuLq/DAqn8u5rk
pE7IR7tR2BdF1dIDtDFH/IJEy/knBbFyRQIhEsD7R4uHkisC1wLyet2kYh9uL9tlgRPXmyE5xdv2
MHNk1KPPo0P3EanPfUsPb3AWu83HydteyvUZGPypz4dVffTfk1oAAVfiFggqQLjpwKxfOtZEJBYU
nV3A5MNbI9XiHSyn/nLDj/43MKRXvv8tmqrRSJJh0TR54i3DhmyRGkw5mCUKrZ3D/UL5mHMc+ydI
yVLRLBpmGAMc8755UOjMw6x8DXpGnTzXHD53KMtItZY/jF19zm2syANqX02gVMQTV9aFc00VZOs9
nzW6ihiEhDe8ZEdH8Vy1MQOPG8MhGio/7kfnongKjt3fSn05fBoCNOCc6nGqgLgy3sx3JdYGfqkD
d2fAvc0Du9OJFOE351r1pgE1gmrvIORa4occOnpmn7ichrVUWh0htPpm438GE9+GT2Aua4SD5eQt
gv9eCNe83xOZcXO+DVJNC6MNVqoTesjESSQcsF+3/3IgnHnsxbfI3tQBH0+wWdMdyRlf8kdjECT3
hezPijDVfKy2itfSsYdexFmjrni1nDqKzWjlhBIvPutZlsIMFjF4LlcRgT0BwNwT63MOVppGX1R4
8VgBNEFpGowF51eHuomCSI8lh1J+AXudwBlU/Yby1UsL/vMUqZQ4jB06vli7fJgrHb+xyMp6f2wk
Lp/8cCGEQQ/2yorLjEjHl/uoymqCQKlAIUSX9JUjZPb2H1AcVTKYwJIrn8oVJm9a5Es40R4bNeGH
lYptBvL1dnsDmrttePfmVJCMPPLMe9hhYMtIFS8oxDJTMf+OdY72r7SWaJ/w8D8hjDP50zll/+ey
E+zwoLTfUYJi0622pkJOM+qBOThzJdf/Z8WSI2VTQreYRKgHXHIJtyT1ufKtVcIDKcbNSGBPjFSt
LqU7Dwn6EYC6TCMz+oR3njhYfQB+KE9wUMinBk7feKtst4gzf7/SCI/mMBT/IRWsFQRN+M0J7Lwi
e7iQbBYOYNzmEZB5NzX7Cguves8Mce0isFHc9hR270rgRs1wfagmSiTmFThT2SDc5cHQ0KBax36B
QaMID/2WHQeXJ2liNP/6JhyT91CsYabWHhKxhAnlDJuEJzKROkKOng/ctLCsId2UzxdX69Y3qUgb
ldK2UkV0HyEkwZqmucCIX5Jgq1MV9fRFyB626Gi2TfJ+O4xWbIOAXSZ79OmHq1p9owxkaouoyZBn
bBQ9H+3N9SsMLBMVJzdDLZRl5liCFt6QvJPM60WFevjMyF8oWQ/BCSPtXsiVo8An5x2d1oLYKmEe
2vqNjoihLqra2Sy504q22dXtExoympUh2ZgPFBrDNxBlz43/9m7dD/cJFPpqsdmHGo0CpuL9WNlj
DdNFCymuuwbIfN+RWgihSqIEJG7RsZqPsHosyULsF1PhFLws9OKy/eVPIaxJzoGwso+4iCsrb/3y
Lt+CCvoTTQFCChV/Q7oVRxfazd011Aws7qlFefJ0VvnLJorTQ671sdzNhn0ZJvKkArKukP/4OAxj
E0S3UfuMfPSqNq8ieh2mtwBmDkcO6231PunrYXvlyxvcj2rlem3QBZqadG5JBSOkwV+dvsmV0n/I
RQyVURG2kIFf0IR+UBYynhGIb73r2Mf7wu7Ti8IR4SMv2AsTfHxdwsShh62IZfLnCTxK4hhQlT8y
hK7cz20FNsd9EmPix1SzKpeVM11Lj5H+deD4cW4cz9HeErmLnG9GNlHJyUM7qoQCeZU9l9GOMeo3
AZYTNsFKTtPtSAo7HnFbJYsJKUjq7jUJOY0Jf8v0iO30i2rRhfscQR7WiCsi6lMW6ctYzlK1NU6+
kZbYQLNFTED19CluSPQmqNTw3U6H97yROxziCpqQxCRJtgKbSPYVkXduYkdwCWYfN7J1zpZejcle
o5Q3kxsp3bMMV5WW7dy3nMt950S5J2DedTEizLItkKqALYMGJRrg9RTgcq80KY3S58jbQuY884Y8
VVD5gfxBnD3qGtA5WIuZeoBRyjslVacQrGfMfs616afG57FnVXUFqQaQ4uHKc6+XI5ikGiiCBi7O
eEIWgzOJYeLUd+nL8hCqQvL1atrEZS6uCbnXUVR4/FbiIv1eflI7riqOSvV/bEgLQecmtxZWu7j4
xM1MVGTbEN0ZdT0UMMV2FR0rA2nbQAWpfttKzC53KcOgTHVAbQiCjl5ZZIUoJzceBSkCDgUGdwsk
C+8vcZCUIkl0BM6Ph/lTjFnG4v1DPOimuRNquu67TGimaT1RQFT4Uyx7qjub8PdW1HPoVcYjZwkA
QwrkTf9UwFUmwZgo3g5unV1qL5cdJf04e0YNwIqER/Xhgt3gc1CzqTQyAEVIKBCmquOLD/yzBogW
B37UF+KJo49YN9MpT3WsKJsFRhX8JacfN4vJikhmQvLgPtcCp3wwQcya1rL9NhXJSYOAUvyNFj18
fnNgRfSX5Izwki03tzIXNALmh/BXytGYB7Xr/hExdVHNCd5mBFfG4D7aOsPJKMmPQF2lSkH5buUd
INv8TZGwfVH7dKqE0R4rPj84Uqy/+/Z7SISs29pYruBFNoQJvKrrke04D8bpeAhRn6ma58xNcW6y
u0OivaKkFOhrUWTTUtBGuHKCq6XJOOtWracFG/TtwJM8NLPiUNV9F73nFlarjdNV2HIlnQWG4w0P
iN0SGy9TvqIXtqzsT6RNcShE2N4NVQn9onIcyC0Q/oko96+CQfXWPf6zu6+HH8Fefu/A/1Qre/Ij
m25J5UMNgg9ydRavRIHYD3V6dOh78nvF5MnIHEJtFJ7spWur+Zac9ykmjkP3K9XyNubCLEfhKsWt
6TW6hCXbKbCY0BclNoWOncrJ/VV5hKM8ovp8V/mLLn+3YW853SIqjy1ZJdjSD0RCEuWe3Gnne5jo
jZhq9qH3tnCuIaYz/7mYb92C+QmctjZgg6F+JfPAIeS1ErRhRQcCa30AY2GUHFyVW3kyuSzEzQg1
1nRc3buclqQvYqpW/vTZcyRgKXho35oKfBtRoCzu1BVXYAggIdLWijLaye+BOOPDSLtGOFlAeet0
GUsQChtF/Nvuqf7HgOV8NO0W+iyePPf6ATL0KfLzGUSniuyDsfziiMz58Porz66Z7m7OFqPytzAx
LUndlObKZ+oPCMm4DP2xvx8up0+8UeFos3x5GeCurfayXce0k02iHqqu343eynFk3MLqDuBTRLZQ
tuw/4hI/QTnIMp+jsbEwRJw+F8dV2yD9P0ODkOkobq49ODBEn96BIpaglQfusE2aPKxv7k2GYhL9
x5fINrec9zSfLYLrHMdOxsRLkQ9ABpQ/IY4Zf1oANW3+HHi2S2eJw39PU2iXPaVC6qL0i5tLnPQT
ckcjfHdlKkWBVcyl9GlIBbm4IGBycUc4PDSnCfdA9Sg2x7GnR/51BOZ4Li88j51YviCGO+sCma64
qhnOCxZwVUADsz66QXkKXQIdP222gF/tyML/vRiBg5olRwPZr0WmJ+SPyzn4YRxcxUocXqf+cRDx
Ht/QcWM8oqRbgsHqqZrpMSUU0h3lEDTqx6TRKXW8uBjz833PSU++JIvr1HKW5IGhkbajvL860jQm
LHr5ZTXQMLtV3ddG8t0zXXlGdsNy6Q4mNHM73NGWw9gtGigXly5Iweiq1ZByDphUTXCxzq14njQ9
IBysO9w5nevgTPSm7nIVrT5hW2DF3mTEYYijGOUgGcV17yDx45wao8GfMOu8Fn4ldKjxBNhyI3yv
aV99iWE2p0n/DS1crfr0+KjvTO41yRYgkhFeHjdJbswl2n8a/EQATHaFgeV1wD5b/tdvNrv9q/fb
VTeYNBWeiHlQ+ZzP2OtY2fU18ULB7If8r0GuO+olbmmx2WI365iR11gGq8SXhhd4DjbM90xYXl7a
fYlZittzzjCbNcJsgSQgttdcJYo6BBXvLYfClMlMKrh5AzwAgImGnBK/wHjGbX0wcYbn09bY2Dj5
VNH4QuZSz/W2Hq3ESnJ3GhRbmYpMOmB/OXXQTmkMFc5uOlcD+SJEFILsB/pp4q5UGaudNF+Dp6nB
JG5wY7JqjYdfNU/AUdNmr3ztnpWSib6P/9MQGu8WqqFNMn3gMmI0eOsX7Axpgc4BNnSDPbyeNxdE
6xgWYut174fNnsbn1+yk9DQDeNoJJp5rX515RQFCiU9FW1M5Svez8bBtCJm0S8VpTbrd0eMDL4wE
flPZLPPfGMIbDP8AfRHDfLEqRCQINC4TwSJ2+p81zE8ap/7qbLb0P7aXS/TLI7i6kvogLTXwqeoB
pcKxolAIsyw2exBsMJggFW8d0H0W/8FdHXT7AuK4KwS6CkL5shVtiPdmGC22oFN7w+q6uGpKmI8+
dyaQRQiETqUmxDSjiVLjeB4E0dm5pETf27BNAVSeuilHZAY3KKGjIclG19Jst1ZwHnzCAHqMntlT
oJN45RsSV7mxxPtTFtIa/DvT7zmzhDnrAPCR7BFD60V9sfHuv3BahdVSgVvS88UeTzG+J/hJjddY
pHDCJ4NOP8YeG9Pn7qe0CL/T+ig4SUttfl2SdGakNqvNGmyaBEnlaDY0N76aI5AWSv+nYFTxmFdD
Wg/GwoeTdRoeouaapBY2R2zqzYSLmehj2XGqNzFEo505BD2W7nX01CGYXbJaJLRfgWVKYSwmazFf
2S0xKYB4kMGBrwhGLDT5wpVzNV2z3K7dSHJBmmHZT+HO56vssV6H6gAS5ZaQW5zjrLZVW+S2Ypwr
bSDDdS0vfrmMcZWdFeFSHqtUk2nnOj8gXdkTemTOOltO0hbrDQti1cCLrPw/zXORyMamaqlgJgZF
bfrf+6EmwVGBRAR7qk/duBg/dF46j78Z3Nd02WfXA/bemvcXWj2U0VMD0fVA6laNSKo/ms5eO/VF
e2EjycYbh9FP1JUO3H1XyAeIVkq5MXZnFGMfsoK6SaPzO1JRK40cUEejDgF6S5D2UTtfiaqlJKdc
zMfjmHxhv6r27Y+6JeMTyENwty2cOHGvFyKvaPvkxeJvC+0DB0LYWBhme24oxH+gLlwFaceP+h7k
edUlYiLadeFrJqeZk+JH1SL9NYVJDZziopSssSXScKK+4qytbdThkmompojq+YTs53D/2qqWU55+
OW619M0dU/ic+hoJNfa2ULGe9vHnlMq/ZeBSj70fHr1CWNt70QqNuS61ppwqlIpWI66FoHxWks1E
73thV9FxbXrfD8T/imi2KBlh01/EuwONTMH+8sFE79MNtYYGKDd15sIzU+jvfZtQKxcornbCuyEx
Z57DMVJR4BCVYBAHZUwZS851UUf5qBsORmCTwJv2Mo66YbOs66f1mpFuZywJVnP5qcjS1pI1rX0k
5MdndKN51DtF13LZbOOCEZnMkkx7JeyhVXnylrzS+fzvUXpCnbpfi/8X1WschungRO740vS/0n1c
vZD37IA+Yhysycrq48raKx3rPqrSJtNudRX+uAwdA2i7H3ZMfkDSf5emzTyf0nBVwbyLYrDY8WDR
RHDIYpEiLe10kTYmJytobgt2kAME758/Me0TPoqfP4gyIat7JTPrONrDK3eWRG0SNnBJNfNV4fP2
nA/J3qT1LQIoeurrXJUN1gHtVMlgouwKy67IsSQDV/QDaB4mq8A8LT1kHVHde3baj8l4Hc+j/v0B
GrmAPB5xhu21GDvLcMF2VJmpgPBxAkigin2DU3+j7q0nMuqRIsOcnxuBleJL7FP3aIngxEXB2myF
PGED0VJbV+NforCVcz4WDgw/gwBX4aYFhXbjcL4x45alw7PB9glPtOEVz31mumhxoN/RdlCptNja
2cR0y6jD1lC4P622FK9CIWnxZe7gaPU30gsG1SjvLssrZ/frVrj+T+MIR4fMcJXij+dERhil6sIZ
AFi4SnIf72WxahHg40FvOVaNALuB1Y8apx3rxLT0un5Zc6UZQwU9596r5BIJN7xylPGilF4/FLsC
NHB3X9GVHnT5DSVX9iLDmYUcL6fKSDY+LUZgtGuxRM1xvFrklmr/qG9Y8wCD+YbUGbMwq3aSihMm
d7EfIcz5cKGL5ZUz/ZxJSzMpswf7P+psbz0o3ikcJHh8jRWJuexurgVlkCaK+B9SGCqh8dNcy3Ko
iLWCug2Zdpjh7YfdTewJNMvLLMEvvWoXOoX3CLkEdBwGckZ5YTwmnGDbbeiHLcIkaPXEnlgUga/v
O5VSxoQ3EBEQA6Z4NR7hD2EY+0wPW6PdWVUCgKacfEnEGW4pF469rOUD1Ua2fCB5s6Ec8p7ZvnvA
UwhtO52BZagInaadgRtEqJT5wwXljmO5dQhxBDBMZRNkO83w0+jCtGnOJWElFZs2Ljx1jAg+FlPt
ZnVv6fUmyoCK9mbE2r1uw/erlMxwuEbZ5TYB4P0laSl2bba/akDliFc7IEmphwT9HsuTIW550leQ
acWPow2K6oRkzMwbbhuhPkl75b8rhwY1sq9/+pBU6WgZXBF9ENuwL/PoGonl4X/L0m365nCeASf3
+/ANay2rvb0XJUaGx5+1GV8AFAWl63PR0Hy15/nzINhEAotj7ZgKbQgO5a3qsbe+52r6zYcZ0jCH
0kjcyUvRuimWXxR5krZJLJvU80BH5QWBz2j6L8ynr2hlS/hUcC2O7M3iUfXCUgSnYb40ubgzD3A/
jUxgIfUIqmNfVOGaj4IcD9riBwy8DF7pacC6g1lHye3/oY+gsOwO+iWnSw6U/QhiZ7snqg06Yr3w
+IhxRsnWDhayRwPDQ0oKil2d6bRkFp4fspmDzn/vv3sLn4DqU1VhCxAShkmYXSl/0hjwbF0jIuIm
GM2VIp8XpdydMSa0ZeTxNsjwQfHC1QgTHX0pOUmoqWHzRp6MfdKYz+ZE2hl2/S4OV7FmGjEF0zRU
H/aOdXr4QTp+L3VR0c6A+ch4z5QCzFM82mTnvyOw67XhyMnqoISdj9WsjbK41jXGzeFRQYzptw5l
HyhQE+xEmgIY8p1cDAKS16BUoEIb4ZZjO3AnZLF92fdE8xg2Wl5xGwy8fHD0Y/86ps7d2Q08m3Ld
SpsPRXSlXLYM1q4gPdf+yv/0OZlPVliHBlVTRV/PjKx60P+8TA3F3hMx7wJ41/0V/IE2nPuAzYDc
7tuPduSnqkryWOZm32QrtaxnZRukVmiJk7d2pTzYR5RP4lXn74/dAhk8BOlWbGl9+rIe4SmWTmpI
dbRUzhNUtuSUIF7rpu5Xhf0eRNKAVc5NbCIx4lpP0rUPN5nfRsCtXRlRrCNKuDIDfLib4jn4/uBG
ps4TTt2TXgRW/krAVDnkKFV0ovjNqVtlbKNotqy1FyqkHfQyGio1KMPSaOHlBzYB4hdKlQHWfai/
kU/OGS9/wARbuQxNUjXBUAwwSenNJcd0HCO6TY2y3gfrvu3n3dTJoLYJZm9pY8/KKR5x6UUIkE2j
4YpITL2b0hSqvhO+V3h1v/JEd3MkzI/CTASOFIcsMV1zctkZEREXPPIYl3VBgfSqrxw+/nK44C6Q
JdCg59INXWG/cgI3fywwTppSMzoZDd7cHsmpQVyJNdjELCq6t1ajDOoaz2gnnNVfnzKPZrMjx/6u
aGZ83PrvzS5Mrtlr9ORxnNQFAtOIpLwTxd7SJYqaBWa3WSvQdbODf2u8Z1C/wxlFmVyhB3Mopb4d
VpV3mbUmgzXbYyG6TlHJo0+yvsSI1OxeSZuP+Lhyme+w7PydnvQ9dbzrkFK5m6wPJ+fiue02p+h0
0gM9FIowiZZTswaa1MdmZ00IV2DorPjk1EKH2lmmSJCtToyf2Rez5ZPiIQDqZfXh4MeNRHfO74j4
oI17eK2S7xNnNL2sSSxBhfmUFVcyTRhOVwdcI+0HYezFS9dL518SMyLwaF7Dpjk2PwTUG4zMWl/k
IFYAzwRaZU64+CZL8fprhFNdUGqOAPpal17MZrA21a4X1WJaYopoe7C6w74t5smXITr4/7vCTB7v
/KGijnTtB7/KFfK4JYYWCF3a+sHMIfmzf9ds7lFG9l41i/nBkl6/M+nWSxXyvw6S7ODQmJllPkwy
KY3iNQQlG1ydxqIW4Y8pdf6aAOz4Ba9oJyFAS93tbuYywwQ4+2tHYUHm/0C5NH3zIqA8aLKnAYQ7
44RdkgS7BxHbXIPvhEbsUnZW80a/5ATMfMWVbStGI/KdQtVn9bp5uTD+vna12fjPmVAIdQbl+YDY
I4jAEvu15FzfRQEzXJSqC7InyVQmmZUTsWP0b6bWkox9lqwSXefsIC1ZqMiRIMqsrV9glXcNLISg
ahayRdN4hZM0u5qm5wv6DSAilhwQzrinLk6W5BOMtIcThH8xqX2VXxX5au7uRvWG137Clq72p7KI
Qnx4bnQBPI6QSS3zNVX9waub3+/Ax0HQAXBxX0y/AmbgF+HqVj0mJWZHPW4IrgmrVBniCjRkd0XW
iCtotigOcaTd6O/h2HrIQufiyyJSyyaIBjRzioFYp78IlVEwYhOP+xoKRk7B5lncoJCVrkZAvQ9M
AtPjiUtF3tENifGYu0f8afLFOXjJ8G4hTunFHAygJZiNvYPTlTo60SJSEWwwTkN8gz8mzWyeJTFb
YRV1JBJWo5zaN1WzChM+VfT/ZvnO3PQfnUuHsDqPVSll4DMupyQwdAK7r7GeKV3gIFneXKv56u8K
NEf+AECMkPhOO5bbqjcgtJqbV1XlcsM5e3Drj9Gqimm8pZGjJD1dBAbF/3LETnP7r1BOYfmM41vi
EhgR0BdQEyumUhdJyhQ6dhMg6hH/fT7SZ7GHrN6Ql9WSKgc8ubeSQz6dL+XQZRnCadL8+d97I5J2
z5uxhV+ESYyF2WyctzrMuiNryUOsE6n7Oz3txGB+BJ6APdIXx9srbITMAfngB6dh2+umZQWJmnmY
vyU1L67ilXd+aUZ1f1WTFK6BPjig8+8TCoiMfacklRxCS1BNn62XaCvnLMUmYeVx4503KWEYL+RJ
KTmQCcZcY7RLmLS9NBnrZLD63NfzhXka+EIsJ7q6V45Q16umxc4ZsFeiqlMQiTFiLg5Ri1ohAQw8
ehQp7XWIpP6qHUpVYhS8X8BTr4GFi4OobE9xQNGpOTDhkHe7R+sZD4avVLbICqyzy5JVMtpZi+bB
yAJQO89O5KrOBO+HCYCGXfFnzK8fYiwmpIQ8bxjrjHymfV9hggmXwCIGdMbYF7oVZ4MEIdzuu3OP
JggkZ5w5sjAvcZTHI+w1A154tTNboguB3XS3BKXlyuXAg1yxRlpRhtnz1sPvEI9jmmTUiDeY3Rjn
56WECjmVx/6yMy36Bg9X8GmwB1AWU4kDqkjCdEv+8ZBR8ZdWRbYeV/05Gy8Ga5No/dM2zQtFR9zm
cu0+tHJ5InBQEwfCTMBuLZvZ6F1wJPYMzKRzBocOEtlR76S+tY/G/ZpDzOvJjaWOPYijENoDySSo
lPaC66Ky40NLa7gH9mxugyWgkyjz6/Gyj0uenb7WOTlwh0VjwjBe8MeDje9xIUSWTEOlC2Jyakvp
YV9fcvmk7Kqwzz3ab1Pi7kv5xPtn61u+w3W6ubyzhoNrpME3aPVMkX7Qp/QKULNQ5a2KmEdwgCaU
RmcjLrSJgtLnkFDLe+Yst7xG6+rMuedRDJWWj8Vui1qphTY967dkhyF3H2/JV9SUrqGwdJlvX3ul
9iQQvfxOIAEU1q2MCz0+tr/dZrlVAVxaGHXm9vTXP2tX09h9re5ym/t2vGxiOJSuyzU0ea9n9uVA
cYdriSMF2MW7IpD7PeTwpKeQnLsEay3q5pGsQqho89vtTCd85xH06Pzww6blIbx4fcUIIgmgProh
wU4U4ZfD6ijDLJcYpacqZQNtApRJZbTrujmj/YN4bHBNjVfsFHAxORqrNhDphm6cGoFRCFkVM1fz
kPKLHUrXQ4EPnG/psjXoqp9ALSZitLjLFF+3KK8PxhYzkdg5mE4LdE0M7NIqxTHrYkTfJcwspVvO
QiefYKSGX77tXxKRTYRkVI1OLUl5dPulsR+1/AIOrlYqn7Yzdf2wj8oZlEod+QH8C0ND79Ycdo1F
v2Sy9WfKy/lFogSK5SAYM+unE7bLq1l2fDJ1jzGf4tcl7rLRulQekYIe+DX72N+xpcaPtmCfCkq8
1n+eNU8IAnfeKEAqMUrLZvcXIOTytOiTUBRa3y3q8DKiooZLw3XagN6liQqMW7Nv6ZR2RlFkDpfr
6g+ic7Vwdtb0ppD3iPYUeaK1VjszrFNjtz3vUHSjm3m8x3YCMApLu0AY6TZsIQ241YpDiUFo9cXR
m6rE+G+ARhgNBz2RdGPyZ4xNmLdoYgbknVJ27Knijne6whxWH3UXiogWtVB20HWZzV1BmE6ZH6Sm
V3HLftLVbkoNH1YDQlR1jWuvZD+nFw5H80TMEp8AJTYE6BsAdSxsbNQ3r1/VIt4tBkzZPM8IsdrR
qyTp5RYdNsiDCYRf9Glw0caIXRzgMekjfWEGcx5UlEfJy5KpsiZhG6wcBguPd3CdshWo3u+dE9YA
ezMLS0zacIedK0QpifwhqRobIZgaLz0gzDfMtypgg8Vv2lf8qdf3EYUDg6jzjbDr7xRtxwVRXPbF
ZNN44KWzGN06Zej23GTa9laVFDg0E0GjwLabRF9C/2o/O81AfaWdDdf1Hvn4gZGFMiONdRoNML10
llhWBw8LG4FYE5GKJQpWu9+z4IwJpEfanRNSSjcX/veUJYTEKuYk5N5a/WLizUn9YzBFZqhA0RB0
XcBa7Tr3AQMlJ4tjCT7iA1r9C3Hilh/ARDHuN3UcWRKvI6GWf3d5oYedqr7Sl1r9/Vdp9pHmynTe
vkp01pqyPFvoDzsFaumnTeX4qHJiazGVg7xW2sJYhyvINEk7RFrxEtpYUleF+JafZo+/kW+gZzMW
2ufyp+CVj/mifDCWESM3tLpliDW6LRszlcRTNGywse6kUffu6z9yHp5f9m3xdNqpuLBKAQyA6KMY
vHdX7abRVKUJVwXjwqh03+6Mrg8wtxNxOzftEhkXkiNExxR+pHqiv4fWAhntXJK7pb43kh35sI8K
LEqW3vxzlC6cx9EqqAtBiUZxb1MPeFYRVyXV55GHyxQZ9bseRXK6CV6+Px2TQMEDNCHrYlWoaGF2
7nmtfqKqkisD8YOyLYkxjaLn5V4hb5OYnziCmKm+I7plksM3vX7+2eAjLWDVevdhCBaNcCvbjo+w
zfZ0T2kWitaeSYucBM68R0aUPfC9G7Vbxhb7jxB0OZYiUaGuNfM3th7ou5jdxtdchullISMHj2tR
nPwA40ojcFDXQy0hQm7v8RlQzumHltDNDZOtDj/aPysmKXCaj7BS84rtsaJmtZq9t0LBMtrr8uiD
sasXjbOpDCDImhN/hmuVBF280KKZ97T/jPyhb39+YR8YCbiaQm+HidebUr4SObdasMZpeVQtH2VM
RYl4d48W1Y2IWdLBAfgR9YqDnqy2ki8r3qq4jAUGJsYfM/55sziQ9vIaRO1kbz/REsDBxK0aY7fs
jCbObqa3JWhowb679I/OIQmg8MXNtDCBk7Q/APu02YjwlaYD1rhXVgEM5wkb6aFb+nBl9jwl4LFx
r1LvbofMjSEfO5zSxmd5KwfgeA6k1blBo9KDPdXEq0hAPFAm/7UcKB9auMbBelkLMId0WdMSrpqE
ZNdDsA4ZtYKw8aDbzj1f5p6S/s9A63AXmMAPd5v5otqRExoxa1ZeVhGZvY21S8IMEUTm4P6ySc5L
XpQmV+1KI6Jfg3eximIWhX7XqZ890eW6KMNtjR4E6jd+aslXCuB+I66FuQPQ6gkPppyqfoEuiYS4
vvL6HkC3ksDkO8q/EmQoNcHauMJ2nkfgbcrfD8gLxBbnbwTnDeSw3n05dlfIkbut9A5LBGj+yhBJ
N8r+t9UeaZXLg6P0cok8elaxU2zXZeHWfSNolFgFIIJIujTIGwRjVQQomjvJIo8HN8lZuYVzlMsd
oxnhwradFVOzFqr8phlwlzsc3c4qIApXVJDmwWm7hEcyMT1YCFBZxDmyO2pNfEpTzXHL4VSalu1o
37n1o4C3ACxTomobMmrK/OYKpznkxkLo8ff9pI/8bV4+AGoXGIHEgRBW8eQPIwdLoj3OfrBBPKog
GrvgLElio80jBudSnVLZ7w+A7UtJwaKm3HIyA1aLnTaRiuz7egyRVYjDatKtr9O72fdKJQUQYvn5
+kk74On9mqTVsWWrv5GvrdnlRjfveE5jNYfFGhTx6taUiF84wL5yAArk0bZ6KgSvx0UBsgFwYBiY
DZUm6D5Jewj4o5E3d/LwHuNJn+opV8toVEQkXNtqbJ6vQjfU5Pt4ZN6MPGLzo3u465TP+JFngUIP
+Sbni6Pwy3eLw8IT3TTsdsHu+8oLIydT1UvSoGaI3Qms8LJcXiHY7KgBjWurR0jJ64Ru537eOGuF
/J/3XPYTlfzQRUuyw5kTukMTpZ2TULqd17YwIZL01IuvPr2Kkkqa0ogeawLm7JBDtzd9f3D+/5ih
P+oXLFCZl2VjIT5ppCwdTZElYmLGs6Ita1RUkbTuCg/ZIXqNViYbdxj82zDwETHdgH5ETgaWVUV+
C1q2dVJT13yKRqycY9yDo4xbfYpcNxI4G7hSPEl9ikI6l/T5Ljksy0kgZibqsSCNHUptnwhwBgr/
IislsQj2ZUt3mxM3mXNlDZW541pwGQWp8AguV9mHy27xJXYUaNH71IkMsciUw5IBqmednBpkP2Zj
moA8S4+F63DE70qKgwvuJd0ENmqJoDnpEKREscc7RiTAAU7pvtiQWl1er09UVYLizdytJ1rKHGuJ
AU+T4myfriaynxiaimSoIJYn8c2vF87vQZytRTYaY46O0mq1aw1Dx3iBW9JxUJ52D0RX40ZdSihP
PUJPGksq0sAnBzpAzSQ08AOrdcIXYLnbzWzsUwHVYCTKfIxABbHci145qSwZCbeSQT0fHjJ9JlSz
zMYSOkth9G5Rwa6f5W6HPYmwTemtKlREIrCsMwM9JOke9O+nAWId4ioYMTBwmMQX5HyTBNpF6c1O
nFah7FxpOwPw37sr98puhtiAavIJgk9JSXt1mku23jM8/e4n6lkInKnaIGMqcq2NWFWWqS1ZzE1+
IDYYwKgxrAvJ40mejSQaCXCdUE7O5EB42zAOdsd7f6+Pct2RYc20hVPlvOjX+iFKJMwTShQjfAu4
A4zsgyVozODU2l8kFwmthKR+qI1xfrTY1/rqwSqomMVypeCvuHWewu3RhFubX5EafbMiwAdQX8kL
HgK8DR+jRrld0Da6smzUvauUORZREMjvUeafjUo8yRWJZ+0ht5e75rQB/nhOHc1YQ8PByaRG8JtJ
CRVXrfkMnsreM2++loCwOfi+RO4FFOMvviYNWaCCDP6IJyrwv07WnUMN6fifrzLU10/tGzwjP6lJ
B12mi3OY0XfwkpYxuWf2FKvErZ5XFER0LsKk1KD3HgjJfUNXIW0gxqy5mEaWGEsGfctROfnihIj7
n0Hpnfv4khdS+uLGAGVfAtGCIXNukSlZ7HJ0aOj/GCRlUhUIgjtmul2IZ/RbBBv14wWPcNWDcosc
KJpyercuEeb9sBP3KIrY4+tnKhj4pm1TIJX5Hy2ATXHLwbucn/z+1S3XuMb7+zCwS17vnJrPqgHc
vQADGUq8kQfVaux/+as5nDjVtXIk3pebEuU1LUzGmbr+AXnyV4thqYQB3n2TFfpxQ4oJaRngk6CL
JyF4NBcC1xyT4k9jKzxWRsejRY3kL25YUIGO5dNkZtKZIxXqNV8DnEsnhHuTssf4TunsEHdt264O
CgaZ1edgtiI66c5A6sWVBr1JikBbgK1MjTfUx+cK2TFiHL5voT7d+4e+Ke8YQcDMkDB0SZdHWm+U
tkrWeoPRwLqbzwOrHcZpxAMp3eWi/EJoqXE8Y/Wu4wbOEYjche79YwHV3toHwb2RU3TL5kiH/1S4
MvfQXoc6LQDpTFJYA6III7YlLMzZBv6xPPIUCpPtyM3TCFNkM/TYatmlpJfTAN350CV4XvSxZv0i
aT8sBko4oYOZaDTIvpRED65YvTO917MOgilNxbv5JR4wC8DQ6o1s+k8y5rWtH/20M2HKkRB/gEw9
j8BloTv9IjKWnpnUayABrdiPMZMYpfHTBc0x5JkmSYPtMcJCuvRFrNAtb5d0E2AHQYx5UeLzibNy
jtjOwIlUexuMfhrRMWmhf6Z1oTSORSWtdMwBYbKHT2BQ5PnG0XHNmkuNYCA/mgD7ZAXiabLS0n6O
4mRPeJNqVnviiMmxgxNO3A4Sk5S09VlP42cPlseqV4ai0EiWzKzlzINPc/FCcgKllpuxvMJT2y1a
/MjjumoQMBgdZUVIqq7chuProE80BPNT9cnJEa3MhUyb0g8HsY3BRuJIxeQFVij1jXx4eB01RTOu
j6dIIUqSbU3qF4qddoe0tekJOwUxnDl6QhE9W7vuFHz+E5VDuHLJsfgzSq7t7N3Wj/AHnyswm2v6
Occ2ThyDCXJsNfeXHkL07EKLZ0azFRRMLGdbwOSvW9v8Y9uTDryllmr8sptZzBmD6kW+1tNX8f3U
jh6cY+UERyszRpmEfJ5hyGSmv6b0YIiMK2v4RXKy17DAcLi+dlEaegfcjt1+hCnBt0zWFB+ILkdy
W+IeQ+kbGqC7xOL8L23zu9zUbTl924Wyd9cqjjHClcI0Jhq41xb5nGFdvMfxVNFwpzV14P9Oj68S
nfucBP/Dp6n+WFynX42XY3TqFtRfYMoiCdQ4xTmzRLqAtbO7stLquT3SEkaMRDurzIyADQYNizeF
sulhu/K2dVA4lIjbUWHUF5O9DBB2ShXYdvPe7ivaQARpWSphBUA7FoSUyrdbgn3ADzmuFiOKJ0S/
8UHk4nULlQuUC71TWvM87AZWP2RSphONKZhAZ2tMwHvfbaELNaB3XaScmHQ0EdHE3V2OFDne+G/F
tJdkTbHNEi9xEvY0lMhdcyauh/1dkkDN6FmHARqe7KM+hTIQHm/REAYU0Wo+RHmlfSvjVjY0Y8Q8
Ys1PUeC4arW/ICYWjmq9i9FdVHMB9zEP9bPE6n07kd4xaGqFBCMXT8H67iR6k9myJvp0qdwpVs5M
IQp0/7hhYR1oASdCFwT01mrdMSTh5pRGTf1oJM0KGLo9jqHbR5kavGj2RWCAg6uo7LUsBtsK++Cb
md/jfx2+uZLqoAKBDYykXCli7WDvcDgkJ3Qqtra/nIUx35ZOPmOD0kOjCXw2mv+O4hfvZUzuKcIW
bbZsxdjH0N3L1y/T7lMYgewszAIGfVWAdSIDd/dx1su+MRey2q2TZj4yQmH8+4ytk5F642xbP9ey
wtKstro+jJKFe9zsygwMAEINgZfuCyD/0HT6EB5LZsjkfJzmfr5izZGHkPV+fYP3JB/4rXfCUL1w
Rs0XgwxdVKvWSSCoGVasNQBN/aeeHdM7XxfLjaZaW+kXqoyn9cHDsr02ObXk9JNI4QR7xChf6VJI
u6JyTpU46Rc/GFnyQklGW2nyhOkS/dHV1tA0hhze4Hk8WsjZH3fTQ8WSq3K3WmWaXpOdmLQdPjUF
weP7mBqsBbE72g5YxY7STiiuFUme+tb1mqL9H9ZDaDRDAdEY9D0wIBnOZ3DGwEFl7NEisrPTNyNt
X1URTXdpGtwcYgm8swPLBI693QnRX3JKchDcCYwTrydzgutwWt19fbjNrVN2J+zA8AGIB4tENzot
aRcNGzVsYC7Te+H7ekurm8iE9JA/RnZMpI+hF8lanXLOGkzNIIOqqGEgP67r4gJx9xL4lf2w8JI3
VWzowc9RPNRNvZ45T32FUm5rySsL5bilqtdGvg0szOlzLv2zMzf3tbsn5EhqRSrnRnMr3X4e6v+R
yU31g0q5FXShsTNV5KcE8agW77vmi0FBxZ1+QEXRNRqq3CMzkWqHChjWRUgke43zmZXbnLSjYJoD
aWlfBx+yMohW4KFuQ17WcRYDMjAF5LguGRgDBmf9Qjbht/4NE8LJknmTq/JrqoKJvVDH5x7sly9H
sULsovEYXT3bRt/97t4ZxCsTX8jbbfdjhElIaSfLjiBdUvYIEAJNk+MlQpaosOX5GRdmf+oOjeHj
Xk4yzABAjR5IYyS0hxOdnSuzoO+exQx7rLjWG+WuUqH4290LziHWenY42C5WWFcDQWtUcurm5r6q
i5+as+3ARaSoicuG1Ip3wKVdA4z6z/uooNzEMtqehteltj3U0HpFkv8Yt+hmMNUpYP5Sag8pMfDK
ozTlZQapo+HnDVCwA4PgpW+cRbdBbaaAz+EPPLjlh3VPFlgCVsFLWVfgF4WiBUR4zsnEoRoXd6oi
4Ighghgfq8aHXk6CwFjSxV7qb4XQVdrghrx2UdlRS80d/XdUxkzz4whfOtVO03sJGzTH4qufRGkO
QJ839JVY38ShqF5n2352rUfL3oFFb9y3bRxf5wcTPJn0jX+K8ifA1vr8KUIljuFCVLg1WDRO1a0A
L2TwtIKr7uPwU6ebTNZMZDjMQ8NM1DHPaTdRm4YHJdgePJFuafif69wxBh9T8aqNKeOCr6VfYTdH
hBnrYgYorO/FKv1A2ta0+xoMCRfMiabINoW05rwmgv1KMbxd3/xILzTgBIhFZhUia+TNtPBtv0cn
BbqEA7P33xIvzt86AHidcVBUUUMezONsPG5kk19YLQu2hxlDb1FYKzmqrgfMW8OBr41mdqdXW4V9
y3JXisZUqMXolTgS2ya3JTFn5e6K9DlPpUKnsyrfGL/0B266OD+1NgDl+eNtAl5DfNOOgrNOJAwY
Deyid7rJ9rAwkFcU/sxpVtqd908z3Yg7ZQ2ri86I0BA9WXxyxjh/ik85qap5mgJek398wC0FULkP
6XDxN92QmTfJHmHfzkLizEdgwHWa9lqRW2fcElkdBSFOVJQuv4GYTBHnF6fcfT7FGrICLzS5VQjY
YBfdwYTFER+hg0JcgIaQaCDMaIc90JtOoz57qTZj5g/vkJl5VEo47meLkODPI40MVO/HJe9gzRFc
ErZcY3uF46AOBJQsYbm/R/BOJpY0PP8jcA0a/kL3Ub2k6xndhNHgdIqLycApG1r2w/A5AQx6lxup
G+m4XFJJ5MaPlghWyqsgbQiO0lbcRWfSnCMmlL4bEUlT6mMlNeOPto5nm1GQJugSttH6YRJA+hPG
CbGd7COfxB+zjuri5sYl7oeUneZ0mMkxbOLZaWh9q1bzTyc/XHLGXV63HOJdyqAN3eXYK7xI9svb
lUWRNqNvEBNMAefFFM7QkvijBJPubMxZ4QwyeDb1KgotWBtgAGYHOAsYvnXxTZuS28N2K1j3pJ4Y
vW/5gFmHlPanLUf/m5mG19jFPBfr1Lqg0Qntp5EhMXhX6/8P63ulJ6z/j1CGgYYoxJsNAniat7aR
HACB8GxVUSURrYXrbQIyZXMf7lNk5/EnHUw17RjD2iZCcZSaFR1/SmEYa74GWKdd3x14sHpF5lEW
7YKSoLDxkLMdmXZeiDscSQr6Pvqmc5w30spYgzluc9NoY/TDwNGV8CdH5VT+kfV5MENdTBReOHn6
ihdYTcG81KtAMxC3YUoYPuOlku/XSsCHX9231/SEypyPYy6eiDMiY1JzptjIBmOMzoSQil56gw6e
xAuwl6ckq1I3FQbfRTxMIyMuCrnw7ESZR46nPB6B2VNkpTT3b6ACQT4dGgw52KjWLzd5+kwQUM9I
ugnhxsuMjNVc7iSMY1enmYlq0u87fbPjTIcyDR2xnn4qypWf4coWDcoi4V5JAD/ANEOapE0sDSBO
+slRSwc3meSJKPTsSWN8JU6ZZen2ZCmZQAbHxOjhWYUH3S/P/F+XhEdWh3Qf1SbxWlP+0/smU+YH
gBOh9t7ZXLWBYN3+kPbvhuK84Sqilg2xXPsmOnl2MZI3853uAt2M/S++QHWPsCe7swLw/Z8NvFtg
cMdFYbQtVqTBCb2awdlhDVKMJ3att0KUWEdaonsN+Y5SL0UzbtCvJXdjII9FvjGfPGKq2h8YYcM5
ydR8WSVfGPTb0P5xqMRPn4WeGHRSLnwBkx6y5u/zLLRHU+6ASVKd47Vfx4fZKrnChqBThUy2f+kS
sO3FZubRKW6wvA45z5H9arTtSFqSE8ZCvuES4iAvaNeExJnOBYWwIZVXG5kB1omIOIMw4862XGlu
gRbGbNKAmNBV4f3LSRMSAho4wNmanlZFjabW/3mNXwsxtiWGaQt7qVtWrP4oOC3rMYBlXHxy22Ga
CHTrBNwbem+S43BGN5eGnR6SG3wCx1QkxSKhDnnQ0M7rRq84+5FxDXVg6y9c3USKAcNqhFc+cuXj
38CXrqyg6NKNdN10w/tABJlfk0YVBNU+d+LTakIoQa9BCWB9YSKYTdPenOfjj0SOTqIIGRNaFOLF
tgfDMscTwZg414b0vzW827AT6yN/tW7J3HMkFAIUaAAzZh6M6o5k5QNfEL7uI4/z0xXJd+/Gc8PV
qIi3ESzTgMWowbqPwJCKMFjogbb+Il9W/peiOJVj2C+nTn7vPOYFuxy/grlUG0KJEpqmssJ/4vhD
I+VkM+b/do4E4S9XdWhsdpIcHPuQzWfEgaE/XNyXr2vxfs/2pqqraesZaoeuTksF+XeZktRxujFk
VnRn6tieFrnUdkphZTevjZBsGO3I/aMsaFmNV3ltkBVbVeAn7xZOkGcmYijJBFuoU5LxO0AY4h/Q
lrqA0jIwtWa0o5oV2E7sPZ+iOkhtyNbHLkQrVtzAg7zB3qgEvHSEFQkJtO3BQ0ejpu58It/fzYIb
JP7ViXgWm3FZKoCAupTvXO2eRmcj6OgkAyTXtpwbbyBdJhIewPFEF75OAZhmDz5jp+M9pNAE0KPY
XyYt5Jy9TaG3ZFHA6hCEtF9raZIk51nytmQqkZpMToJzNbJZAeA7kB8QJ8XyLhzjWSYXuFACaUMm
aybEiDbsx2sObcGKhYADPx7BSGMr1ZUUN/UJxQtzO7/dUoSDrr+3erc4FlzAbvFvXVZRglDXl+bK
QQg+bV8VxJFPe2Aewq28HUzH85EEmhay6Q5msJixw2Gqzo4FPxzszrR8mt36IkqeNWE3/ydEUAzV
m3IqsnfGKpF/keotmvN/XNvPAztCWr4HyT7dbjiSyqiOugl/iPHxNc9NrkPgnYZ04Cq/mo1DoT8A
PW08ZaEP7R1dhT/PqS17K8bd7NlYDpcwRquueYftWUlqQO4sMxvy4MYMVDS+Idwyx/+K0xbo10TQ
h77z5L4uSCUWeWlvsF7YeJyfVPASLfhVCht9TOq4VuY8oBRXDBhgbuPHBVs74EEmfKATlBu4N5ob
khUFEdhY/pYHvEW4/32IVBcCI51ClPaXjVm97//z6TNDxyt5KBrlmAX+M5So8Tyl8sriP2WPRiW5
E04AMmPgceH+VB/vONf3aYXWa9EfsCeTuCiEyqUq8O/pXl4gzB/jVpFBNjNgF0wBUKuMiG5o/rFZ
+w51dOq/UK74HFbPFm0FQRwkQxw6DdJI6lD8AU0GYaoPMO0uzy287p8HrB/7wn1YAj67BKFC/2Ok
2X2W80dXuVonKgzZTZGxgXoAE3ajn9qosDdXhn74teGMJMIC067/PWfh8VRrnPsGZh7NTBiL7prp
H7PMrbaaifCxTrFk3RmUPKB6lfEIbTp2dnhSjTqOTrDffLYU+4C4rP1Z439VE9556BfmTvO4mrej
ET9xVYMn6pSlRQfKT3rpE9d7nTJz+GoyZbfv9T3i5RfiZ9Kbz3n9PUwR2t66LWn1HpwtjR5EcGIu
XQa0SyfY9r6BvylogyyUCvUjXJcUjIraSZUhT3i1agEffbqYMCI9fVF6fVxXeDGjSJt7zOh8W726
xMepTJFEipm5YSh7R6+ICm5mPf3fTdBmbBeMQKKeOGlcAyb6z/pEuiaCtBfB8a4vobV9xgdUJV4e
anisNMLojF09CgI0lSH0n+ElPCzbLrGS0ekOyOLI/kaTiC0QDu2u+ksQCQV/n17G4VKyWkN0EH+h
Vh0ZpLyPYSseUlXKD+CT+QnHJyN6gF1mJwBkRzhmEwid2guridYFrEg/erNzHhjM3kHWIxIKfGhW
pG6t7mqwUWrjPbj5RDjhRWltCmXuRfd7Z4xwhQE+EHEOJFH6TwYrLP9Pt/sddBJ9fwpCoXFkVORM
r+1oE2kYor7FdAI6XUIrqhobRFtlj3vKAx1MixZ9O+ph92LcrhDCRBKwJvrO0ukkHII34N7T9YyX
mUYh4vrqHXjy+Yaxtet8089WEIAnOiox4v8ZgBntiFXoTYopYkAyzErc3DDk2tNkd1lQYVjn3aoC
MdB+W/ozkRS24hJ7fIw/wCNP6fqj3CZxOUvE81wOH1ssbRU/+RXeyKLrWSjHOn5vBJuvE/ZR+g4D
TC3ZhjL7SPECdHVnfJ0ActNeP3vQSfgampdKRxDaVnO3U+hMn3OyEj3fKnSEEzciNw58IHd43SUj
Ka++edHRLXe56MJ0VrsJr6WpG5Sx+UyiTwOaMHDaIQOs4Znuc8ycPDhHmzzK7o8wOxjTUoBbPbBL
yWZbQOBO+e9uQeGz1ubgUubVyjqzjUcR+TkdZpxdllzUxfxNan6hu4lTF88NQAS9RWCNL0+bGzIy
0y5SPTW5TXpMa4eXyUf18IeHGVcTkwByXJOZpSQ5/QMgY5zEbKcr2G2WXjLNOqRJ64Dnel9tuZKn
5n52EG7qpDmCn2/NSWDSK9b6K8llbzgOJmvFNwz72J1x52JBW/uLrVUEvZfXymU8fEKJ8gEQAzOX
djdwPsw2amuA7o9RZS65nt80PCYW3ggwK5hgQHkogkraFmc4ojiL1NmO5MKKuyZF6SXhlwtMcjB1
QGY5AviRBIZpM2NPy5evX3gxVG/jfXwg1supWJ3VPSqRlXRvOEu27AB2MpL7CR1r4XB3FP/z3fVF
QT5OmcRVkhqES+meNNOD7S5PYbKUsXXPorV5bznjQ+l6/2g9KbEmxltN+NDzQIUheMhQUZySO8KE
laBn8Ph+sUjoDPt72f8lBaWcxI5hHO5+bFHihas9sLl6caiPV1/kh8Ilt+a+djaxBzDHZAg7MDsc
tecuDDu59aSl0ZJK7GiYWjqUy+B0JbPjnuJr8ZkIoFmxTy0oZOmSdFoS03eW39TGIxos1bahRAez
eEPKA94CbFUtPlmWpustmI8Hs5MawtD1MSBuu5671cd9m9yf/nvMNxuLSgBRnUh6ntah89GK/vXp
q6vWk+pF04VN54iWkH9f2OiFirNYtZ/R7Tz4TQiGjbCeCwNTZLeDuQY9VA9smoOCzSyQoH2JSL3X
2z4lna5m/0N9IrYNj4wwhR93rm8XRE381oY50+WkTmNuTWQmv+48B+pleVa2SSeMy9M6JCTu/nke
gGuD2dJenUDrub4xcy8SBMv3s0JJC6L6SdOfHTVQNZa/54q5foOxDFegwl95uJYJkmmFO59DpGNW
qormdUisAFkzJLMudopIopf42Q3+vXAhWZpfwEbEpymKtK8jyhz8Ct5o0zcGiMnbQRRu3tDjbnHM
hZCPKaEUNyUBd/V6W5hN7rqlqU/NkgEVJGDR8ILGq6CL1sG7SGw2oEb+JZ6zFHll/DjUWYaF/SHg
OnLY/JEh+vQMNvIcmkewc96QwNg0hEWe12b6g7H3Dahl0di5J81FhoO+EYejwCR+jhTCK4QCQAhp
S/cxEXMAXxP0muCe9rF4wCZbXhAdyk4VzmrxXgohaAJB5vBClEmsjBG0xWsEz7JjVV67IZFYOop7
agIP11Rtc2uh6cPXpRuAsPsVeezcMezb11BbE2Bq6lmoVcj6mKp6V5ahKcYnNYGhqICRCbFEM6O0
f4CWVEa4RQMI00cWvF8b+Q8RAYUC1qfCShxScwpVekzYmQl8kIo84yHAjL/itGmsJ7QvJENEOu3u
9FHz3OgajRDTowOjftJ2lZq03+hQ7++LWGtmZfwney0ERhvoLkKiSlohHWgp4/r2zp+nahm4JrXP
LAEdlqWJA7gGgvQ5DxF5zfrOrxSZ9ykKNBl094yWVrVNZ9ScKxZOsTxiMW/K2QWFCtuGbt3KHLk5
V2ztJHRl8vszl6pV/mTNzPsQsxe1W54ALye8GmVjN2TA1QaItiuMsUQk/g3wI54/c45mEHV01B1E
0+y5hL7A/huCSXtlFGpr4dlRCeSgqKOWq9nl2yPryLKHgVKtd3JRov+cWDiTFxRHmnoS7WW8d7Y+
c+DLgKd8KIsZFFuiW97B2Q7KCYIFi2UhGk43mOYUQ7pOnQJk5eYPh8MQRJ3ewjM5CTLRvOoLnDiF
U2mLOAEPWzHh864+P9ctkNHDddNAxmpF3hqy/LMUa8uSYgONsPeJTNtOaLaFPm7nzPDqCb7s/yrm
22VwyyrGRhLS/VS3MGifBwFmaJjjOHQuSMCFFP4MQswBG61dAysyC5ydCt+QDYnMYEaHbZZK1vjv
EkKoJYmypNB9+7+dxjPJfS0aaMWv+cqn7RwDcjgmVXhYAAFK/kJJlVZSnuMlLw0kDvF3LR7KabA0
OmXdzub4WOxYHKaM2f6AaEtZ/QuPyz8IcAJN97lXHIAKlNeZeCfOzQMLGhYAYVY7pyh/iP2SFfPg
+n5Qzp3pioCmrHTC0579XJX8qV3WXMAcNT40Yz1QQ5oume05thSZkORS9DP6SJDyHU3tCSPVJRmD
3gKzB4PTKpPy7NzZndEbzqA5UV2XZdhK7iH2oZWs/0nw7+Ns29JMoeat+XGXF4I4clNjG1OiwIJM
OzJOYcL1Hb7Wt9kDKJfO0OE2CL13/5Zp06Livq4lXkapodVAbWjwNxlN0NV8hk+yXJKaVF86yqH+
+sh7+ptJCAxVneoJ5LW0GJAP+NNyqAicuvgkjcm0vj4/eThkLkjticJsJo9y1sOowL94CFkENlMk
DWnYlaCGrZFiA1jQIztGTw1T2LXPOWKAmlNnh2H7zdrU14Jta6BzBEkct+rulVtXX9OEjjJ4gpc/
hv5XfGoHAMBDh9rgFRcFNrGJLl2RyQQE+C4Tbo/cbuTOyVWfRBDN3zhtsGsMFBLjcvQ0VUiF3Snk
P/VlnDVpIPzhMxK01rnO75ILB062+cALg+MnvOImWdhdDHUN1Koeh2CL29viJA+AdGwU5dPDEXK2
wDtIFg7YHEnx1CYqI1cUQ4ehpGdPaC9MqRkNkIz/CXEgQy7gbJEQ52GdK2MZprZomjxc3nFtGlYF
8TZpMs7oaU4MrcYEgC3/wzZR2N3dz8nM9KA1UWDsp94d4vwvYgKAwAe8qKsqepefM5KDtiWPCGu4
nqPANTe80KDiSjNUj8RSNzonh8+LDOY4YCJnCwde02Me+yQ0ePi2tjaQQzFo6EiCD7TiB0tYIAXv
hd3dum8UtQH6qeX0aLTH3D9UIvUm5WymxJomJrzqgSTOd7eckGD++8xYxPzv62B5/2BayAHre5SA
VGHRo25jw4ElwQOmt8SR46L5aHvBpN7S8WzIrt9UtOQCZx4tiO80sWG8aAppoTQauVltHgsrQ9ff
s/f7vQecLucVFt6oFastIOD3BkYja+nBOsePyRe0WqqRZo6Mi/No3qd9AnYfPo2As1Eeq8WApHud
3eDAk+hpIldnaq0x1r6V3VKd17TIxoejrDlfTsxKEw8U87iq5rdGWrydXlyh0LOctCNrW2kODOK1
hdxW26H9Vmqh3nhiZY4IgXSWBHmg5ClNVxoR/3VEv0IS+VG5a5qmkGQzMwzgCrrhjPqKKK7ar8g+
CtHPf/+DeJI4hjKm7nf9npd+URT9atfFswcRpPEm2dpn0hMIG0ylaD6gVTX7PzeY/vYSucnNlkJ1
u23oAJvzGxyEwtpxc+kxx9TQrD4tQLcFEQveJWfsZWfimmiopDOmaZjIN29yLxjXc0C2fGd7VkrX
b6R4XYaARoBhSaoOEE2Tz5rBFaWM48byDNh7OIYK8fifyS81jiCJw/d/jEr7aWXf/Ma+eDjsiErj
JWMS7V2hS1UTCu/PRWqsyQB9YOnJdLhFXdR0pMDInHRhi4XV+MGP7Quc93HJlbCflQnsf7kNc4uw
L3uOBoPZpHTlzCr9smfR1bNE390fYFhn9GditgzrfGmK3aEt5kUbPoSJIQabQMX0nBqE7NwD0bT2
QTvbfmqEn5FkgJnd8oUf4uJ9DCtoFG3uMVH5tJxTk9r7eeVMZ8gqbLGKTUNB/pfNYtUZB/WlmV0Y
JSZ3ksl5o27t6piFUPVGBwTwiViV8/MNLE21I16Ted5FusM8uNDj8rWGvBa7wpDYWgGMP1I6t2nS
6rYw6aS6qJjCxfsK/AphJ4IrVlgVXIOG17Gt5mXOR9vAWYywNZYNXTVwHEn40yszHWVDo4LtbJWC
PlOXOyHCgDDQSO8EyDtKDeyjtCBZ/+x2Nl18VuqJYiRvnw4B7s/kIlQqsEyjAVHaO4Tdiu3TYGhi
QOXtMg8s8oud26muyhMFoD2m/p0gcE8+HNG1+RnC+A57nQ7wzer5YAveol94P4avXf06iGGT00J+
WW4g//sPLsIVNDLO8f1oAIHJTLU5qgedrsy4ZcXp4vcXG5B/AqUuejpdxuYXk8MJoVcDBbN9WZRE
VDJrnVFR1+hfi0zVw0cgPPPxZfnwlEYL6HRrASoYB2Vye5jgaEhc9u2ZKs7DTORybMn3Palakuuh
0iNNpwH+Hmnecurwd6wIMwKKQ9lsB0cxXLApQ4zGZJ2DsewaTvOhUQCBuPVzhkrnxPyZ2PQQ3C5P
k4IIKcOj2+I4I+c6Lj3H13mdB+72ZqYf7DvDYcARBjlQtWEmYTsOwTZv+cGQoTLDcnA2iEkvXWWd
9Bq2+dhBCp0cTUnL8laZNjNuBzfQrPQPfrFT372sfXkz74KXLrknJGx8UcVN3btePTP0jl9TD5aH
O1siBcvGh7aIWakd2FxIwTJls7eXnuaKi4yhbm81LrCuzkC6DDJMD3MWHpvCj0Ejyh5f0+GUEzN+
BXOOW+OpoXMjMGXqrAsYY6uYCJ50wzxKxTcsWguuyaWBnXMYP79sK3a+pp+nAROdAb2OvxbNtKUA
G3scdxGfZDVCkXb2q9O5dixXYHcgVO+djOf9RHA75HWGWt2zBqNXteyezx6KVG+b1inA0IZE4jb8
8tunQeZDjhUh3zM30esbSspUBwrg+GUY1v4QfrZcArq8OnJPjmAFVegUbUFSxVtDb+vTxjo6DcbY
2cTomnaDsj17eKSjPMGLnLkOzrlNETw662TTsR/mPaoLV0GhBbpwNVT8Uh0f1P2YBkxKmLnuJgg1
daTF5Ei+oPj907Lnwph1UAhYWtmF5QLzUVu57DmY1rqIQ1vTPHteXump94M+5LaIY+IyNHlk6FsJ
hGLcH9QdQZbIG/4Od5caZO8biOBEf7u2wTSj3tziBxJqMFM+PFJWFKzGGrHQ0HHOtlP5y+2JGbhJ
1dXVkqM6D7pLBdPHsDC6+VokR1MChH2SHzsUFp8Z0SEbNwiaK5bDA9ElX7VmPv2Yhm5WTQwrd2Jb
M0rHks/rJmHjb6P18PyY7ze4mH8fAJodSx9gA9SO4ebHkCv0rgKuj+OnnORX+iwLAqq8N6wRW7lx
hBoz6WvqkQGtiQOSuwyV2GjkQJ9zkjtvkjFyJLIqdCz/5r7CnFWTSZf09dNbcbr5C25BgbzQEr+M
FWwf9b/JINbrwroRV12m5L7RW0Pl9gbMVwenMwOU/FqbqM/hRtTMlaPD2Hr0feavEVRl1lfxaECj
ffAwk0pdFQD40nJ89B0b4NvXq5WUBEckCf4lbm6w6hFzEeTDrQbpvC9yZzEminUdoQxyVvb3wbKj
7M9B/pjczf/OUfNxoFKJRb5rLfnUsk0SSXVgJNcuEv6bvOuaIbYT3zBmO8ChV2jeVu4fycXfXYZI
CNPY7RYAjzGqkBWUYAqYGs/48dJX2MvwlRGcf7sHHvhdvN1Sr2jPGjuNukCFnu+9Yb8K5iZqsmYJ
QK34qZpq4a2C2ZMs3MOawLp2JZNuJeq9QCHjALg5i8U0pYu2FzPdBudDqLgMS5SmhdX7csbM+v20
cN6b4YeJtQME8oU26ehzksVOqNroKIQ8dWqOl/tkGg8Ps2+xBPbX7TLY90aUEhwi+mC9YV4SHPTU
g/I22V7UDyLmXmVgux4qQ/1+y8YP766nJYU5RCjWIuXJXLVuU8IfyQLWhJwCeUsSU3vREXHV+kxq
0h1NDz0bkaxjUemD09H2hO/Na2VEfqIxNMvx60EJ4alR1PlgMyzVzHRzCZ4b23RH2aDS+HoIQXvZ
6hGsSvtAB3oICtcXDVPMGlyXI6ZGgs8+ueFaXZsxmuqxdTZQogwLX/nhmfQkpjvSiBBPjmVBy8Mv
oyD/KtjNH+fKCOx0opYn0mjD4vU0v0Ry0nucsgY9rRX+HDCGpdsSOkawUTMoQoaoYiY1EetAs09z
tbb+naLxkfxt2IQj1qibv+geBgfpV841tc00k83JXdFN0v3oNnZegbFEm0JLpzkfhOfwBLyao6Cm
oZaQynSVFtL0nKst9SlU6F5AnJx1UU68TaOHQ9WGpIxG51GJ/ag21w6ZvDDVdR5AdmULMmLS08vK
rSk4ERXPEe2d1N5RKga6C0xzFVIHm82GbTWTFiHDCPLgfeUG1wPOAZo2OUUhx1TNA07AHUxZCum2
b26wTyePw9b/yumBhy4i58oznbmeSC49X3jfVsFgPV/WYGyLOmzHFJX1fuc9D6HlBBCo7MEcsQMf
SOTJp1oJbsmClEyNq+L8N/psgHWK/yHECkGprY9h/6taUbWXCglaZzFP4jM/vfBjaN1ntVNaFlOZ
mYBhNwNBy28BrgL+y7v7P5IYPWZReulW1fkJlPCvzvBo+EMuUFv2aNLb9EBYA0Pl2qUcFtaGfctP
r1dflUu6R6dq6iWCpa0uWfW03KqA4dsqOADX1j4XLXCsdZfXv/+HgYilmQwKmjCPVbgG4lgrjnLE
szuZmp2vZgPcsS5kFOifOcJYnFBrK0cBz2lb2lesQJJZZSsMs5RoYxHWVSxpfO5sfP+DOxgjPMeU
9CouUI7hw8waUOcamz+mgN++WCgAS1+GVW75r5Y/SD/Pu/zzN2pmlhWdX+e7QniuqDHy3bU6sIGw
0Hycl6IATcUa8e9Ev3QHjvDPOgEWpDrxFGFgPjQn3geIHmbfhCJlobJ/L9wgT1hvPlwIeiWzCKFm
NiGvF/SUCiSd47W8SyAQ8hyx1QH7gg/yvHWhddAbJqcHJhKqw5gjGo7wx0qmkBB0VJBnafKgxi64
PrTGrf6AM1z7kt0wAOA0oxS+u0Fx0+qvvGF8fLvtvM7BahWLBrJSjCoFkrFujLtMFT3EITpNVWkj
6RsMGdWPeRuIYsJhZi92vB8+xatNEAKRRQShu1iilzEILP3koUlfDMWjxjp0fukJ5fx3pRKmkeqK
jXcg08q/Yc8jybUnfWma1KUpZjN9Ze0t1WudViTHFoGazsb2nHV9OwdiCMcY4S7N8opCQZCsjxkg
cmGgFZ4TMPluPC+cUYlxwtjszwZA+jpH84OJU15Udfp7d5i60T6FzPJ/u9Sc5seGZBcPzP/IB3wk
ZKMejyuwo9mnaQOM4hN3p3WbGfOij2qZzc9ylfHizAYF/wlkB2voVZMsEtmOlq4N+DpfX/m29Eu7
z6E7ux6M6mJp0cmxd+zRRifIyM07xiBKxJ4a3dSv1+ILKnAdAF4SGdbM28sygk2dyqvSzolSLhbw
SNZLZUwZHRR1x+ixi3cUZOFO6MOQCil7GnW8HoiWix+J8PX/5KGY9Y63wh1+IsYBaBUzXWpIgvXL
aie6e8Xo+bT3WxIrV3lFmtLk1pdwV//1WnOkx4z0sYRUbdjBsa0Ezb1KTmI29cmW3mDQv0YGeGwt
YdOXG7pnhb/awWAHRU/09DS0y8CIXRXu0mIou1/OJ3VkgDvfKDyVn6aaFxBjYAMR5+odz5gajOaB
KGtCfcIKc/PVhDg8fwSScRO4J4tgdyqPuLqvHtkaUKYd/gkB0P3ggehke2kUokb2+JJCNS7lYtap
JlnfESPdYN5nI3pjhVrYCwPNW7xPbMAO5DfLdWXHQpTkWUQNeQC9gyulodJAWQQin6kfVIQKxEDr
KjGshILK9OWI45Un0uGtAUCB42GwQn9mvxX0b10Gv1lj21KQ4gfMNTxnf1/OD5IvC17jHwNNr/f3
lZ7aUANr6b+js0sW3RE5+CtUzOzIBsDMUHdEeXBORB8CBo1AodDtTDZRMQqy3hZQXEvjGBuQGBpQ
Wl6kNxm+IQ6AywkbEpsNrNFfEn60UwrTI8CyOw5V4F2kgYYhNC+EmBh80LsgVKagoWf9TmOQkNHu
nz8nPLRhbDLqHetKtuYx9z63SRdHcoOJWB1QnteTLGDGE9iMVIN18hLNT9B4R8+UG9PEjrFxjX4K
1r558ylEncW2ilrH+j0ahYNcze0WDZ1/7f5CeTex1tWUHkpitwCHocrHK8W6DxUgo71iEXXj15Ir
ZJQn90Wf3xff2GzuUdjmmjL2YeXLnWMS639wR/ebGmYDKi52GfM1bkCNJe9AEymXioKJy5rvlDZB
TNpFbIyiwin/2BtTVTSPHoMVtXyvEgEPKu3cl/Gibw1dEQ4zf9OM39dDsZJ0VoGh/N4HstOvIxAr
1C+P+BUmX8QBvE9h6x/oGtl5aQ7MwVJUcjydXN8RCeQiBGxyBcX6Pc9geVgwCkpXJAhk6bG3/13a
FvT0Fxk603HhCUmas2iXK0xHtqGTIIbLnzJa6qQezIZWEDfq7mbh0KsvyjUy0bpk+Z/69Zh99aAz
qMk+1wzdHqDk5+/2ErDaupZQxLplPqdk2pVOkYi3ruiCZSw4k95Bh9FMMN1GPxJnlp4UOXG+qquW
w7NMOLB0F4SYAlqwMVlv/cQgui//aoDGE+RHYz5Yw6ST9W9P6tW2VFFpaD3dyk4I4CWOPQ33vX6d
ZDhsNxmQm9KddG5v8QCW80IP7hxabwci4uPW7PeBPCdSAUgzZbEC071aF8jq6jBDRrv919YZNGZ3
op7dG8Z7THvgzXWe9u1ERRsrlOhnF6NK87t91L1gJruRwtIsYR+qqR3GMUoVwCqXM98yB2OQTk5T
c4m7T33sTv3Nyzb6g1jaqyAqdH7fyL27vj0oDn0biR4ZTO2zK/ObWyfTzID+3Y8Y7df9fv1X09ns
kMbzcXTe6VuPFbiF9/Ydpw3xZUDo5N/N5YardmgTkJeJi/9wvHYVnX38IDIU36w0jqSNM8aHGxyq
VQC1RjzjNE9t4ot+CbUBYdqcVObAytpHl8VKFNozTcRcUNDBLU8mjBmqEvMmudQJorb4M2mjcSeG
nvQvBl4MZSWxrT9u/NCDCY4G9BLr6Fb6Q6MlohhFkQ0Yi43swio2dNb7kuaz9IhlBc4lrq/irVkQ
DuDBZekJ6SLozt/ESF30MG8ZA1BhXLhmnAu4XZ6GaDDpU1JRW/mLsVZSQLeNnCDP3LrOmedv259Q
niVqAPmCGyRNk08zFhzJg0a7+fG9mPN0W3uQX5NF3AYciGQYjnrtUMlotNPcz0lTRo0ztap2oA0X
M86X6+xfNW4s2UqQF1VWLgCLfHqJ41PKIOdTqPDgW8s0T/LnepBkVCiD5DAP+Qt+SHqwdvUPgoTz
Tw7feMIaD74RJtSkquSS/+XU/DNooTA01ufT8eja63mjFp1sIwE5wze5orE4r2NAjIwvhbJ3qehU
qLL8Rhkea4gRlq/LSw3MRkwtRb0vjjs93HFP397taTRLl10sUnssJAvMaDxSj6i3XnQLIxeuiYV6
adjIItuBvlDg42aRWSk8h0OrUfVBHnHwgPZPp7i6/jfQQoEmzeI6izF4DCjQVMqzShR0NgpJ5JLT
sE9NK6kO6gKtvr8g5s1Ka/ew4foIh4VNktv8GJaO05jSK3tDi3QN/x9LHig/YuaUDjIG1YQgy9IM
sJ3tcOIgn6RlnTn9ErbmMZVsV52sUv/YJa7/5OvIf1T5E3rmqYCfImXtdFQK9hmhMGyrMvi+wetn
blpgSwiHQitmzVlGBfNBTIdftobXn7pCryvZKOJQ7fxdXQWRZSbUmr7ZRBCed27KbAhP5lAe8cN3
SmSO7YLWAAulxvEbl+LwmiayLEiAdPR4y3ugeYkzeIWucLQeyA5G53ivGBjhzAJREQ5nmZArOAtK
8DsbbtYGqOauDYpnLCHI3As+RAGB7fvZQtUCSWZoTTGIqcOap2gTVy2fGVbCkf3+fH/AQR2EgIxi
DWchwdjuqU2SbiI8oXooXTtFecv30GFa5479aFBQXDqOVhtL8SSLufZlepXERG1qTDxdc7zLkWIp
VKIXbhKwtv9aiZLTUkZjPyPtYB6zzrl1d2tYb2g/dIbvYyt7j6eDNrNNafbtb0ElhtPEcrqSw9EA
7QvIH8uYhxSP4iWiF/z1Btj5MkkURX2c1yBKpvS4uCZoDJkMwEFDrRHHcPWP6CBZ+FRaI9vY6NX7
SeMqpS+JD1ekD0NqfQB5bt2LdtwKkLznEtMtxCC5UkKPNktxP0W7+UKZDWHjKILtxwE4HaSF1iFs
dl32vTCAZaXQypxPqzFg//YDj/Q/xXF+ZJv48ykGL/vi/FE4Bh0zfUxQPqMviGGLNyexx0QjI52H
AD+Fsg5h+b+MWaFcSFtDidCEYzbhj+ytJgaRJVZc5XGasNriyt+/rqqBVUbDTetj/dpsF6ui3H3P
+nXyvTDxP9oRIRuKP0/Fh7aU6NgHXwDJFDCTCcWH8sWCM7dBynAjTIfQNZ6VMhbRNQ21pa2TQaFJ
cPtLmyexnE0/ChvT4L/vIe2DM92yWy+p672gApAqvHN6KQUkmTOkVjbuSaFfEgGPyR6GeDaMcWKj
j4D8NReDr2VX8adq6U8gNIogVPNHsa8BVVal1xh/pwRVE0RgyFdp7C1Abu0uuEzb3sifX0q9jguk
UWFBjFfZQKrK/ESyb4rUnJ+jITi0DJVuCFen60qpH8+86uQhcr6ulZYBx/SehQU9c6dqJm1WI/WH
4aI7+nf47/6CkrtEUmMeJZnZgS0qvDhCCtM4owBZaoOVt4iC+X2+Ds5UcYb7t1ib6swpYY31K7Ae
lPmIMrqWKmSP5SBml0Z679LuuG8H2gWep3GjGXSEzkimo5R+igBkN4yfibyAeF2KtVtGxhLYHj1M
tUqpSbsTVVfaQ0ZZa8J8FGxO+4jxqe2uubWrPzvGFHMSElPF8+YtgTMS1Oc/E+KmbfrPuDi0csK5
phXlMIzk+qQVJX/eFilJvb0mrvW/XoIoGhvFyhrb+WVgwSpwkdhC/zcAMMhJNdlkMolWZ5aKk7O2
F/NyGi7a4OJTLHxW4shfJo8W+5bc/0asUkBJaSPTvevULK6Q+deMDjRy9gEv92ry2hdLVKxeL/eS
QhcpZanPzXRVuEeGUUAuwYB5c9hhWZq1rmNaWKBOTdJABwcvHQUMFd07xbMOfA+DZITZmyhu+pjE
X09/gnOrKxj9Wlk6tfNshLGw6VD2hMOKcTX092sVnpYgdwBKkLQA1mQXF+kzCp9J8MHY424bWbNa
6DxbltX+BaplxdJT0q3qb81Hobq5WMwjZldO73Yh7R4xw8/kQEOc9v/PDJ/7A9zpE6SBUTS8ezR2
/cH2xXaxOYE2uvb73hGZAylxO7RxCj3NpzdVWkeaUiG1tC1RZktaT2/HVjMF47BsBRrHSW8LIpaH
nznKzvtS1QR8+/0j7c7W5DOpht4CHVfOFSUVUJkVsClS8q5Ow1lO69iVKwiwTYXyVrYQ3HKwBZaP
bNbOanio1R7YTi8tcsB5SvEebK/us+TdUhmWUi5v9AtXRVrn8bRLZkRDAhzXKUP6H8FSMu1vefb7
7X1JnNOCiH32e80uPxXf1d2cL0Was86DcarBIcRnH7InPoAzc/2AbxMDpTf//RHjNM1MRYHHpOA/
HaCpN4bI2dsRO8lMjK+B+7S6l0M+x5pnXLBFD6S55Z/Np0rKSPKCfIkEAJgbKYouHwXBErlKgEf+
8d2kgr3VOhn3zaHfXsbBoKqqiyQDNAzuIyQWmpP9JpZhxSL8ZlqcEh9J5DO1DXpb78H39ut6kEJA
6aGpFULgAfvOn3CyUGuoy3D9DerYW53c7ndrQQ6tQvUozOpe4aCLVii5OKJquzg1866WXNdsnBAI
/rVKfcU1PQqn2nKSwdCft3F0GcKfaApACQ0F6KPt2RzX270otpK76xDtXvQh5kv0NVv7u8zgaBWB
8zCgaxOsYZVjaeqp5w+sUpCfPLWMTuwit98goSNDK6SWK/lzqnKEgkE+E3upfw97tnqDkuAYAO0x
gFcOJlBXpxGSqewSwn5L8eapni3MY7XyHvdQJgU3YVvI9EyENLDa3YtqYhy6KXyBixXaxUMz3jKZ
g8ri2MGxMKbWumPBUoEuwoiRJRgJZN+Q2o929+F20mVphqrau5muKM9bTwTb0r2w4bgAfi8cXROt
J4XJ8eZBbI0qzofeCpU077Mk+i0a4rxa5GHgXtnkPGoRwETlSnKt37DjXP0/SxVHYrcZa9eHj4v6
l0668yOrwfKiORk6NRmZDwqlZLxJH9YhCFkObgtOCfmNZuYd9PJndDBWDSk3vRV8DHD3QjpyhW3R
RhDCJuC0l7ZZFw8NzpHJMjIUyj7JuPh/EbvAk6r1JBgfvBwHJ7sJhKAjqj7L9yfgJmV/Y99lps6S
rz5Ptptnqc/HXbL5iYA79FU/rVomcuWvYyK19ubOD0VZsrjeMOOxbxdbdkBPX1u8aXOtrd98E0bQ
SBTGpGCV/Zm4JEbCeb+PT7lVrO3RXQcA0f17pXDJCLuVx3KXmTjxMFC0vEeUq6k9Lf3ty3yg6La9
GJfV8OCTnStBU0HpHyZjf56BAadTBnRs9UYZxINuHkSUN/aL2pqXm2iNOFkyITGKe38hmxSarqz9
eJuJW/9GQ5g4l+bA19kNsQIwcWP0oxmpCk1gGjLMXrhFtEtAEzkPcZILBLUCW3E1AFimF/HUbm50
2XcWVmspM2Fllc7HgA0wMN+JIVsyVVvjyt/B6cP9KoaLyE+JaXoD/GuB8FiHof2/zQCYZej6RkmT
w5mdUGphOWH6+/WzQ/8CItEy+Djw3qcSqvE5LW6sxnzGNh6tyAtDTm3b5FS/epr4W8xAS0oGhhVG
Q3k0bx60GPnf1LTY0Gv0LFUanr0cUVw68QPNtSqzHwYiUit36m0q5BucDil5Tfu1HHuoZ2Nqod1Q
m8roZxoTNaXTrRF7CmaXF7d1rI6RaQGq0vsRBKrsbdneUIM68pY+ZYD1lrn1NSBOgjdvAjsz7hO0
XYbDUycIrif5QU0obhlZltGCOWUTh4FpEXJLls1KhOWLEwFJSelyhq+WybqfEEEKrAMSyn34wBfb
nZvNdZFpB4Ducj9wlRcSBs0cZUFxlt6GC6OZr7fgXJOy4mimdVD4HdhWHP+3AObt1VxtkPlTua9c
AwIPXDJM4CllzdxTVSo6ahKYRdd1tXuhHxBf78MC6HIqwxscQqkSs4mMWizgzRb9R6RKQNRSBaxB
JG81DxZIZmbiW/I68AKDnkYeO01muYMz5QfSI2JWboOXUyIDxawApw+MIjJuu2QszUavY0z/p3Y3
frabAzm/jiV/Gk/r9bMIlViFT6tKi5V/FEB+xm6UszBfrC6i4ZbYToARu7hiuSzZrBYAlidYgg2Q
GaJNptMk8qIGYb5WUJthyWb566dYOqX9HRateqQyWemnTZPvw1W8RBoKtGiSlDxufmw+EoYG6VO9
eYFeA7LScPMiejJzfAmwSqCpAwI5WjGBc5YM8BILbHdsHoUntWu6sVYIiImfcTUjUm6+8ZUdIvgj
EEBodfXMMnPmmPs3ADz6CuCkIHVjsExzvoRCEESPzeU1g9SBT0yY1yjd4NGPPNH1DrDamZyP7KTP
menT9QeeUa5KxXg8zXl9aHyK7g8lM1TVEWz5LL3Th4+yfRyXcZP/o0TgD/Hrh3BPB99mIlXCTdW7
wLvlSiMSb/2DNPevfMIXy330Pj0TCvQHqTDqDtnhFXuyLbd67cBLcdtiOF22dzA17eAA+W7ov182
+LOtFyWlCKTyrAdS9X5/luFRwMFFqHjIiDeWW53Hh8EaOiU+XuxRp5/X6XzP1VTRvK+yYJTbKZue
KxtpGfTTYXLfGIkUTXBQOENWzzy505yZILy4t8OotigTYd2GAVkOA0pl/DY3dkmFTbO3YbyBkcox
DmBxSMNrvDPErxSLneJtH2jiSNscl6NggoVQ8ZGq0ON5rV69HC0LA8HAqgdliipHXCdSC0Orr6IG
FXdD6KlpeiPv90bI6ZajcQh8etL/qK+m9HspbWYc0EPJDVZyJo6Iv+ylH2nP4zkWF5dH+5463BSf
mSd+qbZsxoIM++odMMmDfIKrjERU2KsBU6uO2cuCcCR5DFCHttJguS1wJFQ7xjudDSi+OkbjiwkK
wIPhORcZEVCJyJMcmcFyudXmnHguE02sGi2MZYQ3vWaBSdCTPDnY2t8wsH32rAL+xKBhaV+qpYJj
iZnkVLe/95y5KtFcDpmN/9xut63EEAlitklhajWYk4K8IlBq+9ng0Qv5sjxXlJ3XmzI5Z9VgGIma
YirsRbTUVNfZCfoRWabto4cTFDJyrcv0EBZBSmNhEQevfp2AhVbLAArbDJ7HDW/TzZIorSfwhkao
Dsvc93IXOyp99/qNjuap/obsdbEAe5PqrLTkd9EuoCocGvksRLhth7uU/+r53bMokKp4buAHxEJl
b75usnY/z6RYaMHQA23OmXB90PthVGL5YGpFls7i8vUzroJpN12gOfrh2k4gnv7aZZjlcZRIfKeO
tZnqFYgfiLk0JiI+yrufwO7TxzyhcmeihMjVY9CMyrl2up4WhIM3TPlMrOsVTlTmBgCNJdlk9ZLW
0uJKSWi0k6x/mtMytW4ZlnylI7lpiu4pEav5ludoOWyGtLTj1BbcSQ9iUUJxl32EMKtZkQEkqRJE
22JbhmbjZEq9JSBkVCO5kVmLZ+8FylmbOQc1AMOW9DiB6qgWeoQHPqfng/6L6LVZx3XNELpluDUa
v97gGExpUvXdtZbzfkS2bX5M4xfbNxfhd+fUvFV5G1lRMa/BUBQbU6XjUg2PA9rWKp7XEHunOhr6
/+olE9mgzQ5hXb6OW/26icaGVeNl6qjbckpk9dsxjP4SJKJqUCpRyDhM+4Xin4FvzTDOKP+Mgtjf
vJFExAtcWtkTlCHEhd7KORTD4VF49zddZcZeyFh9Js/0NGJh+x2l5kHnwvf2KJex8PbWfNpKgorH
+6O3RAQyDnTRLnf7ruEWn0zakae66v+2WUd2Ox9yw7cwlGcqLE5+7wGffdMNmlG+p58iqP9w1tXa
ISOiBE72Qtb14VUBJ5aDDrq1LOHg3as69qDWWJsK4y2ObWOfEzl5g9NJbGAXlX++wyE2yk0lL8+N
AeSh4mVEV+lX4ZlDeUZTBRMDYURNp1oiPbDVyZRKYsyxGFPq0n6IBURcf6vawUfHDhGtL3QRh3kO
UV1Z6Q5XZqK95ulHgdLLSYgBS2EJhMWpVJMhVGFoEe3Y+AcKJgoOBN5u0rlRasjVYLD9mqLgY7D5
R8E+nNGnmozQQ1VdOp4BYQxu9dO4Xev7EIp0TQsm+jAwi7oz1aLbAdNs476gFGZ8yzgkZ2t8on+0
KDaWmDGdLPE/QQ8yi59eJTf9F1wBLwtfbtvJUSpQb8S+EULrOZhXlLXk/cxqRS0V/L3A65wkotWL
UujrVz+7aKjRnfFqn+dK7i89pbaT2nV30wKKpHvYIG4f1XYKGbMPoTu9Ic9e1ZIQrRzVnye5pDf/
WcCuR4dDTaclB2YJOEqUx+1OJaW4/3NX4QaPnDUbPcvEA5dzWqAHzJ6dmtOJB8h4xGcGLibkMQWV
p0hQRfNfQjQ4ji5fO+B7oy89Pv5RD2/1vECEjbD9LY6xY2tth3VsPPEjb9ECc4sHmzxUN159Px1j
8xOiZGd8jG4RSDI/jsqU4ihKND+5dUH38TgxvFRjBVHUx2wN+GNQt0VgsFaYza0MgKoRghIlQyuo
G9kK5SvGkiGMLhn15oJRe81srAhsUWnRTIL+Gdl0B5nkm4gwHPwsJ2mg058E/scffuxE/E68o87C
hAv+gSk18TZIA81v8QlmoBsG+G5tFzFCSVuTWHgjTRPZyzJHVOCkax9u2PUdE1f7NVEoN13D5+As
4HDAhbwWfSO7RDg8QJDEAtRLe5clqpx/2BfK49TLxT4MzWc/vEFlYv+xFuhuBOp/MuqISIfoVQl1
6StvfmHkDe/ODO9Ra9rh7PQmHBdB/160nf80PlOsFdiUPjgVgv+YkKM6Iy2znI7NOMDL1E9LYtCm
fl5c3xgFBmGtLsVnaAY4GVD77A7BqvfLZnACZSAiVV3NTU83fqr3PZG7QPUceTg92PvAnoVhEz+g
umm0zZWwog3lLZcyIqALymF+O1L9Qt7VowROcqT+2NjTMgllc1ltti0ShyHu1gAILXVQwPuPp4Bq
vB7VAOmB1jparqvZZ5v6AR5AhAAYgrv1u2jUGjxrOFwlmHt1qP4HEWz+9izTj71o/sYlGd8pEocE
emp1ANqwrTQLjAeNMW6qsL2FNzXQr+VCCriMijYuI8DA7tosMKAmtpeI/9v99MjJbNnKrgKE6VdW
k4FbdEhhMAmH6io0TXsudScSr2onFdps41+AW3cYyx5tDQXu3DMHnlN2PSpn8RL3GaFS76Rn4mxX
rN6Km+e8K/Wjk6JbMScRDFEyMnll9TeCcU+mq00jpmdkKnTjNG+B3l335YF3FAWktnaQWilyeCPE
HC0HCOvzaRFru5R0J2fONHQ9ojHqBFzQqfnUKJ2kagS3UYu/mRPyNjGN/5t/d3JR8vZusRJwIBeO
Gdu3rlFLyluXLqH3vxa64dYHmQY+jfWAeCW57ErXYJxyGJ8d50NRpMnjFflsGJpFg9EHohVml896
UZhhjVP1bS+ev3fxgWO4VDVYCOsQ6yRZrbfAlLVIX8AQlmZ8zi9+GgvXHEsOl4QGwUVEjeNDLHxN
xwUjw0CaovRrpAMnq/HpGkjnVv0qU90NXpYz+ye8x0FhqN57gknTZ8ovRRivjcwho5ygxpW+ZIbP
cK4p/FREfUQw4MXuy+9MitOPk9sl+8kiWhAQrUnHKzKXcZpRnyIIw6fOjqBSe4/9678SU4riZuwU
D0RhUJQHL1+/2bIScfmcBLbRS/U8VaXiP78gIiXtJ4Y+mX4dNA6gmIZUuBB+P1xZAtlhQF8k1T3W
WqDFzLNlgWXP09nHerxoXHZDxA+GBl5TOdzM0p7BQGXODK/CNLJpgOPf0aT7d6QgXGSNq5RT1lBb
Tt4WOLJLuCoYCR4dCTwARb2ae86iamAyGxyt3Kwsl4JRP1S0d7X5olQozomZz/9+7gLK06q/dk9p
cjVuef8c9WIfmtqWnN7jlyJEubiKneGFJS3wX6V4XZXT+io8h1amujzom1/83+Cb6VjU1CFtstzh
vRxCIQ4m5G3TKJysNQQc0EEQuGSh5VKdFv94gwRJedNlL6CGorcos950cxHTVV/KqcK3sDaqLM0Y
a7XlLYtzJnUvSykI608IIF7cdR1BgnyNjFqj0Pa/6rKZXfbfp9lNsXGq7+O8EvRjGUSlOCcg/ehs
/D6SvZPhnsxXeWsQQTc1kHw0+s1Pr5fvN3vMdXl1YqGEzQGzXVeed0y6gmokaz9bn9mtPXz1FQ31
EyDZx7E8LBZKP45ceiCMpqtxS7VrPV9E1yjHIDxDtusbHTyfIgFEp/n6LMHp9vYzLbeo3cpbKAKk
UOZh5E7xiVvb7G9p/5HsckLKtXpBu6Tn6lOoJvyskpDH0utB6rf0dugbWP8IsT2Tfx+70K4MKpV2
/gzzmN7MbWF9qn+f85Vrwx78p2jHOUwEKQXui+1VgKqaur5/In2urCdIUvuwAAJOBaBjtV3jHKxD
NmF0lvl12Ql++LssJ0A2zNvBVDGusJynjHuIJFzkl+/TccnOEjGEWJZVBnGJFMgy3iso539fz96L
OaHi3TYJo9lbXC0UWbNGWgWlc/nPIiH/6OPYqhI2yufwaTAnNe3xSo4uCDSwnNFTKTPYwUNwCKC6
Sq+jXdR8GEN7MyK56vhVQeUhjCdqlRThPjeXMynGFkPEIBvLoFumkce0zFZSi6E40Rb8cafQu4Rc
rXatsfnV2/2VexSvI5XCyNx2YjQHDtI5/5xFmv78H55y9RI0RHvcplDIvcF2XpDtrE/HlpSE0Z40
HFSyo9yV4VRVBsj10DTXg2yRIjNskagEJ6Xs/N7iDbPSK7l9B2jmxjMGdQ4ChnnBd32zyvGNkYME
WVxZJlJvTrY16DjuFeSz7xEykdMnl07ilGavCajyXaQbBgXgKls6IgVKeiUEkNZkX/+hMMIS2aKj
oiD9PaDys3JYrR8T7y7qf9N7kboAwY15ZTsvNRmDu4gDoloHQu2ICwvJX5GdOXs35KxQDp6NET7/
iguNA3JjyPgt3BFCrgbSDiD5mcjwg4522vN+9kGD9ZhbshsnGxkB2Hjzyr2wiNXIoo4o2LkZxvj3
e+0C4DI6jGRu9q7t9prstMWsokaFTueJozAc4cln3PbIcL2KgL70ftqRyu2Z4M2wQ8NWBCbfQfYh
3wLz+P3WlSto31+DBffRVIQReOt/lsQGsoe7Cp9V58rehlge1IJ/se4gJxuBJ143XBQ+skpxdzP4
jNrd7wAHyQlgzUimDWsAomAvHKRyn8jofPcNOuNWueM7y3fnuGfm/EJvyV4R4anQKtiKAiN9p9gP
ov7EAfMvvjBgXKbAggMYCxJImPxMiD3u7IMuEfmX/ZcoilVCi1HqcEyG+ThvI3u+w444ZSO2cVPC
wNkqh0W4J0G7t0iSwXPo2MSpkb1VM4hFcn9UikHq7cTSU19peMy6FIIYBnN7eKctpYBz6YIwj97L
M4isOz8bhBzBq0wrCnm0xVJnVdLgbO2MrutNBA57mZpYp3khOxxOs25Zx92++QZNwnjfopVYvfu6
QJVehfEilrq3XdWC8XzOoetKSAIlejcTrOOIOQ4KFS44/Kp2Ry4jU6fmMq4x/SKOfURVnsT6zvDp
xa7Cj4enHismQb4BwlBJxBao5qhUVJXzAxKR57BAzJ3Bk/rfjc9YUeP2oai1xyACDcy1HACox3Aj
lf1s9YvzWdQ12Kv47W3PZA+TWSxwf+7H/9P+qetW0mj6r7waCPyAlZrUR6WAoWBfvqRDnoNHTNBn
7G8JQn3p8b+UjIEe9tEb+QC65lEDrlv4vKTTF/F5v9Fp3xYmtjYI5Y21Haeu6fII7ehuqmrSJm6V
hN3+kBgh/MyBF7neRKfddaRDX6hyyRfd/tcJMzGnFSJB1lPPnQoU22MhjE4jKZ+ExaE2Ggv2vqC9
Sz+Ei87q0zNal30prI1O0IbNZokSQdsnZMORbnUR5SJBMoss6bQTmyXU4h6flrf3ORkdLQCr+qBg
E2wXYyEZlMwfKv+RWrT1fR2HFQtRqqlrJ2wnhvycQZQc/Dn3A2av99KIiUVn6DiSoxCNW7xelsEd
aZlWXOAMU7ldHmmwZElmJvC7b98+NXvl//R0MFetmvb3VBIIuYuFKgavUzwKCmWPDZYHYfHj0Plu
sP+nsm9VjaipT9xauhcC7TYl/wIuDuPk3/Tk0sHAlG0vQrGx7bQ7vvLG5XpluYATLl1lF9dl170Z
QHT5kZ4Hmu4wK0Uu5Iq5h8Cj9nx3dXkLdAdBhNzbw74j9rAXkOhPnJRYXC3pWYSPMFXakLh04mTy
BVPgZZtLrUOXApXt0wJVnuoG15F3RsAlnskP3gnaz6ExpiH/oKGBWsMsZ2n5C42jHbFK64S1NcXc
44Chgpt5r0VD+pJMcJIUa+zSgzSc240PZDEdfX5TRY0cIklURe+6ZQsvvW0xnN/nJuC/1kZCLRnI
Ij4X1pO+VElJDLp20F9Y+r+XeE912y5UabaQA1Rt7RVllZx6MFBLs7+cReQJtuPZwccWwyeMQi3m
d3Oy4b0Yatbh5v6oLqERt1LEJqEhAJm9mV1qjBpMm7iY40Yks2C86nQbV0GBPSivu5d9ak5l6stZ
JfEuZKcsrmPEtmyMBz7OROD0Ud7e7u5SmGjSpqULygh8YpvO9N/KzqmzCfQDO/RbecxfsZV2z5Wj
gR2gLU0QzAojHOdwct0Sa/Ci/Cc4UNO+TFVaF6kxCBB+4kHNUU/lWnMN3zOWJoFZ8IIxFGrsesay
+DV6fy1YryfmlhA33fGvSItzfYZTLMcWohnl1G/X2ocCB7SYhX9UwVYHIdjlu5JAA6QEp7tcHr0s
9KG675hmi3G0kAskrvdjRfDoJ2DJHfGz2Yn0PyR6GzXD4QoJDsDPEUTfzI30G15yd1l/r8GHqkX0
6/hunE1nUnE3ObVvU9Dc01HPPc+K7K1gvxvfz2yvvj1+l38CclOHVg5vtNdc4bKKnyu455BBC4KU
yTF6Fw7CQCKSi3pqg7GDvSIqZxYrPCffg3mC+i/Rj8P7sdEKeWwWAL9FVvDA8fS2Wqyad+CwlOIV
5O1K2WWzB2bvJmtVC0zeg1fswnubIgJjbDRuZhajRkG7x3iBYZZ12bVtWDbQ2Y6XG2XEkEUuRpjB
DsJu1BHGTCMUQEJ7FzlRVVrym/c3pZHQZRaciUN4YPYet3+wE23hKsry9LEJJiKZl+PmlMGZuYOQ
SxcEHZLmQKcOjwJVC6mwiqIb9DSPvrHxV7EhZif0vsVcfZeh9iCyiu842MMDtFtIfv6rFV5NeEA9
UDYirU4DaPN9PqwyOeLdnJpNpdJPtkXmOHV/6R+WhxTtSCPaFmv3cdc7DExDsC9Y29IC0OV2YJ6h
Awfe7JUou4HSMizaN33JZcxgZRveyNDRPqUJq6nCTOvB5xDv5qky1QyBhnwbfwfGdwo5A/pFg3bM
5jOf5Wt9XwvJBvgxiPoTW8bTXmzGHX8vwMIDqKDsB+DlPIoZWOcqWWH8doaHPGhExyP9QqZju3uF
uiMHwjV7HTiRl03MTSeqQW0ASH1Wu0TK+1xrIt43DwVlhD5ca3yg/9XCewSsq/ojaV7DayKt9MJF
r/12m2DXBfR8vGF/XtsdPbMKDfUR/wLMKfazXHrlVkIERiTy3VyXpG8US6+naPzuRHG8hu45lLqH
APPs42oFXE1gs57Y3g/fykGUxDfIpbjddRdgkxs66KXvG7v/5/YjrpWqEiipBkroW/WBPQ6B376+
UNfwvdQsw3wpuyWL+LC/XMPyJIRZcXCg8na1EfI1orFlPX4I3Vmx8I4SQttL2hX7apQD9Fd5IeMF
Do1GmuiCVbnBjI84r+IDAj67IPZW9K+T7FNBGeq/Wz1ZEi3TOMpicJjoSynN6WmCcfi+ea4Yp/v6
fMQIWlEqO7nGY9U5vAxB+p3mv0VRcQKcJBVfKZSgVsBpadNA0iaNEQPfNYXC9Xu5gpr2DaEc5a/8
8DhCwyK9fTY8M4cLb1co7Qrs8KCuYsVmhwCOl7MqkSMHuFeZc7qaxJRjaAjwPjGMDSMzlqoq1gjO
7rH2DN4swnVhpiCA9OvvQeOIzNtXCT+tPdpSgRwOYz/kKTPZlOoXLhQTlSW99TzdueJK1cmdKvdw
7YEwErX2ePcOq+ckUcyRS9mTwl4FdfxOjAbwNWPC0PHZsEvoSKIBXSO26JlxoRnyJpZXR637TT/n
RGU27A8WhJnRv7ghRrggfCOzDdbmm+32JPwWj17dpctzhua4MyB3efmeEiUr8QEEIWBTCbOK+TaX
sfJwKftCunzxrHP88xSgg+I3wNNQVS7A/PBIr2BjlkD66+VV7eepOTDkwdLrHVQcjq2+x8rVMImP
v15pqPI2+E3Xm7IAIHj2FBlB9QHiGBViun1853deUfF8NoUmQQe4v3b7uPrNsbh5XUEA7ivsiKde
c986w4z8aMGoWssKrJIFINq7Y8QM0/s0ru2UUxprp/I9dWYkl7Q2YXh3RD9O+JRha56J6NsGRR5V
vVP9iT7+Jnx2nAj3/xZw1jWDnoIGH8e029bET89MejcegHmA2WUQ1wf3ZriUev7LSQNrhKkAUxx9
f7QVY3bjnsT800U9BE3BU4lj7Hu8JPphQSVcCqDDBYwd7ez12fKoIiYZuUNf2QNTCdCh5tzI7dDU
IMqitLyF89kRG1OV6AaaG9aA02BEaN9WYYAYQ1zTAsN+l4VJRHdJYd2wEG1tG06U/s8X2fIDWR8b
WPNFH9KyiMZnYOsMpqo90IpQEFc41ec6Yl6i7W4EedRYsM84ysTbSfqLYVn2qsa3xbPHj/JXHmcv
f64nmZa0+inbk8oSauNPsM8rxQXCErrd89zsQPNz81AsSseeAuXhD79bCN93+5Kf++LZGQT4EFNs
kTBKdeIaVmKE6jGChOr/VVdwgR+VPiKcEz5d7QK9R7RPUr/2CpjXC2G0eByvO3HbAnRZ+SIyB9KS
Z0/YW0ZIP8tQlmAzxi/4lET8WYroMqAgYcyDpBxR/KUNq2n3Btq1v2ovRMdaPfRvpxYFFNmAwwgN
GPYFt2g1dl+kCG7S4yVNRD9clXRzazqSOQ9HwLZ7V3Dl+aE9eHlS+a2Y1WWs0M8T2AV6B7iMCGVU
7s3njcXnWJL9STzw8n1RCnrHVUb/7Fit766KzhoQxVvaNCFuGPy4XiOACn6YAtLzJ3WUGPqEQpkK
GMnrlcRKLCh4FkhFyBh4DAfEfOv8nThhyYWKQc/YQyyos6pkNhxlGiiWpPeuErQ9PCypcP79Izva
P1ilD7mHGcc8tnNaAkxU4lF87WJWWaNn7fnMYK6cne1hps+HhdmS3VqkGOfAuvmgJz7+J25bSLoz
0Vtj5u+fgkvqthcH63iIIBfi8fMDgtxQXyOTfCmz4lFw6aCiqGRlF1W0WTJcF6vSkD8b0u2HP08l
365rHE4VhvZC0mcHB28ukHbNDbJ6Hsh8uGKCrPl1VYsobtIj9KxaOH/Cuov8lfF/TUdi4V3M2Jfq
LDrSqjdK9KSB7xofydufEbFHIflrKZdyUsEzqo81A+gFqiSRQxCmooFJAL0bAkwA6+c0FZGzAxWf
TUldnyZx2VGrV0WskZCdFnx8rai0z8L6+hkdK2KI90MhjkYr53/RWrRWYqtTBysrKjFoolEM2y58
K+jgS4XOsz7RVeg9Fd9iMT37IdAbRyta5XibpV/37YIBQWe4rD848+dR1ncFnxtrO/4c9N+ffeQg
CMclA+dCtCCq04/tCnULV58mfeCZJY5+VXDSDSkjhfY7PXdohgrOzQeV0znX0FSLctet76n2cQII
DZpM1b/vSHEFd0WGmGcl9wwInncELxZWqCc6agLsIFQqKTQWdjgr5yJwVYJVd0RI950UGOWIuZbT
DIutQ5Bwyj8WQLDOD0amnIMq+8Rb/T20xDCig5U3MZhFb8ZAuTrmCgmjNmwBlrjjGzpEIuAmFXLK
2Kinpd3VLcGwFK8zNgvkokVmwaaqCVxEHqYLMdD/uh1LbyzBghJq4F1sFZEKyqLfDjO0flFSzdB5
geMtEk6+X3lBzvsVSLjWdDmdb+hH9xMwysenuzTkWB3BwRNNW1cNOojTtvaco5DPb7G7oXZt8Kb8
V0FydrFzZGZOWzBzYhCtage9G0uXYA2ptEIAdBLlWrbMiWA+XDJPo5U7Xb/KDdIoQ0O4as5HfiPX
kWd3Nsssv9GTb+znLI/k2fHyLoPI7Pov7YUa31s+R+5c0LNc8Dl1XIta8upfTOiRN+jtX+xv65F0
8wXWsMzCp9IBlk/41dZP0FZNUOrnBGRDmJbGmfPNQxvKlQZiwL+IZgNAoRr5iS27PDxlElYuU/kV
nSqlPnkvPtkdtoZaekUxtHN7DKkJp4TA1U/hMrgzRlb7pnq1L9Y4tgEx+BLryhJhNfXIkP5Oc3/7
fVjGUCVJGCe66iBBv/4g59rO+/O5N8wAM4rz1d/QUsJWhkB+IYNs3xLgQccpMhk0pYVXZiDcFrBm
Jt56Rdqca5RKiU8qGlNYVl7b920Lx5XfmMkEWt5zj3vp3lpV898pX8aBZsE3SHX0zjcpCBQuf7wb
ExJKaO6ShcCxcptt8lWdekb1sUmfieFTS9c8Pkhfve6ERsN/tFm5RM5VZaCTz21l0CoD9tLPVU9f
8bqA1gqoyJS2iczQDPqmrhcZOj8YlDScos+Xu1uIY5VA8ggFp4bbIFyyaqzAZnxaTeJPuGVV+5Vt
L9LV9+7ADHqTc16cvkOvX6PSxb7aQCbWh/dcF2wnBC2k5Cb/DuUwXSmcGXTMihNQfVVPnlWm+NWZ
yb/HBfxZHiR5nfbrqObGKP+997kdAoAJR4nic82odeEzFGrk60F9gO8rsNslm1/irNgjnMv26mrv
YjEWpOzgFPpmnPKBoomBGKsEJ/MX7f/hkVRjMKYmEobkiHNA4XVkBzWyU0dcf241V0aDy1YcSmmu
WWBs9ma69Eb1j2nphZudttf7FCb/6aPn6MIWS8c9Qe7c3ZJu49U5I/K70+jjreRioXPF0XpyKmGv
t9PUtLgGS2BTPLZwQAh42IdHbfks112OBlEmPum1jYYl57NEb7kDhPVj9FWGFjY/BGvNtHTvayAM
XPMx6y8sdxAcR9AUpP7+9QT/fFSnCfDFkARjlvCHHp3SYkgxvorxzjNB1kRQwNg2ni2YZioDzeQg
6OukD+OmjRGHVjgxQYyR38xHmYV+XZ8pHgSIPLXBuNZPi4AARoyMIxCcPwLFo1LbAKjdeX/QK9Qc
ekBoprPWxpINycMo62jXeS8pVFRdtkbe0nFtZ5OH2AYahz+tLzJ5SdadFzyckYw7r+NkABsTCDb8
9cM9AaTQcXSAi38M4meEOZczwcgDpZyPCcLTkwP8Jn4TEP2wa0WuSr6lsReyxOWjEHvSw+iHCXoy
HGay75Tsf83Hw5j48UNmYvfZnnAcjWJHtlOqFjrz02AOWSoJz+q8ycbhdBFDLawZWJHWdGSeQKoo
jElDttUdZz9zqyKi+NLMIirPpUsmTIYzE2thg41n1vlGLqgBV7kwiTgQ1+8mdL+ITsVXkLJQLaXF
VnIEMfiQUmI5ppBmN85VdVOtAVf0QSIv1dr6oQQPz3bI1hFXdMFSkDO9PrWJVQfE9GuGnBYqIoFW
fGOdG05CEw0y/i8qufTd7fDtJSU/M/Utx+qZFtsIBp0kfnVl+w/3vf6BNuBzZm3uvdRjukDyWHqv
cE+hvU4Y1wG2/3hzoc+zi8OmtfRyXSdap9XFm8z1iFLb9P8UoVrzrB/lZyylSZ1cbtX8oji5Au48
o29rKUT1J7qgKiDM94yCapOdalqhT4rZyAq8LLlU6URdinuUANDbhCWXL4TPvbmppSaps5vmnVjr
WgS9zqExu5YA6a2+tjH5xhaOiO2VrFBhQm2kVWk6Bs1oAtlmbwIoM4jgwqH6RweqP1QrFWRXwBxV
YpryNaj0tyEnt2JJwGtldp5Gg+ZLSeBzaDSi2ySflvwpuGep/sQNji/LSD43+33ZI6gTu8uq8Jl7
MGQevTzEW17d7t0u1+zh3gkrtZFWUTbMfnYSnkMDpQyU1JH8GfWnQ7MzMCk7CKSR5bY3v7DdlJUK
+iA/u2GdHnaWu1ZU2HyYp0wVXeKLvoYHB2uHLFKyarP2g2mQoYHeAKtR2kuYXBeZ/YgTzqf28Y0I
hqU83VnUxavXTFPnvW5C1y7Mtwl/ZvHxqViiM07DDK0ZfLX9N6vTMqWbUgbzbx5Qbs7pk287yVEC
wz+pW4ILrmbvDXeYdmz8ZqfyNkIjApZVexX+Vn9FT2sa0RnSQkdZ09MgdMWEkHouICeD9VkTywAA
kTk8Ovf6Q+f/YYZM4s9fe/w2YW6gkqTNUDKJMnwG5Kin5DLIrJJfB0ZO+GWlhG/6MUhkx+qZrb4R
O5Jq3rVISuYKM5A1sLwwNNDnHcTz1pSFtC7Vx9V6d3nkPCrcjtUFEgOk8nk6g541+ZDMZtj69WqK
gd5SSU0fQRmphp5H/f3YYHIW206cWF9j8fR8OXE5wwvwaL8INNWO2kGIQe9/pXC726BC1c2OrHjE
t/5nqZEc3purqjJSFe6rpbxMJGMqsQBzrSY8t5BTpYtpTkdxBRaWFpFkrjVZioNwJokJEXQAgrQj
YKzw9XbLlXTtXRlqMxDXptZJkoXQ8rNMGzuaxkroiYalm5+S2Ud4sTTjIoW19lsIC1VQodljUqG2
gAxS3p0JEGcilOtYV26H//BGKJmTuXdKp2Fvxuwkq7ETetVtR0OEeYBo5vSgL1iqUgjCsZGaL1cD
r9f8jmLaY+j8fjrzjCZ62rFId4pyPRBXHIrB29kVj+ZvdDOIva/lpo3nzPJQ0J+v6BcCw/BiGzBk
8z1jqfrUzV/uWM+RwoIQrNBCjmkGs9SPd4EH9hlTEDWFAOCjYOMA6jwHAiFHBuAF5AIETgroqIAQ
30G452Gwj5daIca/GK2bN6HYQKdJOpYf3Y+Miu2LArXgr+/TuffqdcMae3DEe8YXD5PebG5wMVVQ
cm1yy8SutY0GbiBZU/BybIAtEpHJmaC1EJ+oX8IvGG0W4dCZL9uCuhof6ibKgKMiy/BqWzkuCVov
bu6dRd/lR67eVkC/dSHeV8/MI1zck7IbSnE7Vho23/95WNJCxhELMg4CvnU3SHJWyne+OkCKg+QI
JbjNBgJu/2IAlPIjjm1u2WNdReiKm8WQWm5uQk3bipogAWxkAimZna8xdsXIRJUYVQVcuBPoEDtP
+PjcHovZMBkQPbG+goZkl2JP/LEA06Q6q3Iov631JCCGkBDiKXMUC7DmpY3oHatIokC6aj6rIGyE
FjVU2uUxx04Hzp3mIxwY6TUFeJrn3NIxCboP2TGlDHCJSAe0F4QK0319mNjKtuCf1UPCTGHxgglv
EREDjID2+xGivIT0fsEtXU2gO8sEfn9snXBcm2Edz+59GgumH4kv0/MA/RwtTfDRYKsRVgoImCQm
eH0fb5TlDGwT5I2fG6EIAX4Qd70SVyzvrrlREgMNcOeQfY19n8BNCyX2IqHAueHeJIYmm53a++kw
JLUJvff/cYkfj2eVyQr5pvn/vSos7t6S7axTrG97ylE4PawQHjFatVCifFYAtE7CpKVwPplSZpUQ
5SiSctvhP+rn6fE3L9If5U5SrDb8xer/B1lZ/22OWVv751uYdyWEz5mIvvW8z4nQKTN6jtDTMcV5
taWJqbltewOBNlETqIDyFY1nMVRZkJzTR2AxLMyFKQOP0+5oeObbTTL/1JHEr7bfZfNe4mpBCEAJ
4YW71m56AHMY5TzFSLFLm82v0bCgdGW5J4pUgsYTjXsOo+V04CJl4AcfH5JG8+7mq+jlGsw4DvAn
dD4uQsl/IUUXrOUbnp1CzQgESsbbAz3vsNZvjGm00AmgCjHWMjFlCx1wXLp5f+FjMSQh9QdZ5uUq
mLM5TbAqCLvMygzAIsccqNlKYgZ6hOx6CopvjToCuKLlWLOox4RHRD+/bC6Ldi1yNsPdB6JSVbEq
G71D0P36Gr4mDvfKzELDOFQQvmR6J8ut3YuhUUjq6ALzIKzwE7sIrWo5O8VZEMY6PfCck8EEJOtI
VAPDLHv+3uGMWLEkhyivmZ7vQ6X9aUepTAdM7/AXEdWwLymoPl6PTTEGug6hkpK5ryeNiKvfCd1z
l55VYZ9I6L9WiXfH2lCa0qNSfSASnVBh+8+VINl/nFpLVLwsGSgEqahLeKdtqPs4QXKyUBaYmabD
45FbfzBXxLP3uQ5XiD6jjgQ/B9URX8QkcSqaOwpproW0eT3RrK1QfTubuOlwcSoEYNb+iLXQNm4f
UD3T46SBLU/U+sJH64OAv6t7XW3lnKgGJu41RZe7ooDgeaqkPeQcFkb87/Aa6hAA8fzrg7LiHndZ
L2GjUn3lSZ6IL3CbA7LZo9BztoHIqa0Omwr+01xUJHBrHoCVaz+u+1AQdOG35Tmcfx0v8QvgqI3o
sswDU6oG3xlL5ZMQ+5Ft/9Uuh4B3QjolS6Cb34NV8/Uz56QIey4cr+8/XaGl1Ny1tlcIbdqQ/tSA
PeIMt2oRwkUpufVvXAwyP3Y3mPvrZ52eKoC68mTa9xcFWUx3c+Rils7aJ6tNzki/87TNWKzSjpLm
UrmH4YiZPXLcvvMEFdOdyUpMg7j0Y95HacTy6KmKjgHvOLaIH4kkNlYRDZT1LZyG4A1yq3YO/Cxc
T9KGsYdlf9ZhL8WhheWWygcEfJmMHOvrqtW3HHIKeoKAqLjY7UiwOelmBq7hLIuNBrMvNwagLcDl
hrQkrRS0URp2AD/GmvBGUZVGsFsFJ7mMUV3RiFIVX1wJhAnHmix2i6sldxXfu7qBvrNI79Sv2Csg
12vsrWKfqI9ASHwPw8JDL2eVMs0dLQTagib+r56oXyJcMEfgAyhiCH2mNB5H/9DkwETjMQncX48U
UPPRGPOUPhLLgaCqFaX7swdTygrmAn2Lv4vg0mfn89WPKUozXXO9NPnOtNKYoYDKKz+y5KIO8K7h
SG+WPH2XDqN3L6OtHa8Z13SnCu5cU1hm8I7JyAMDtLY+1cTmKqvZI4KmvoIh5NKu4toqgKuHYiJj
f1KGTaOa7JPF326UjKnYZ6SqUe2TQdDhCxFTSSbbDJjbk1RqofZKVhvRX2+dAGRgLoIwlDUvZ5zX
2B0P5plaYTzcQAhy0lkiaDmWqkEl/bSm/OYduR6S3kf1pnbkeOdhRgeywb8slm8bvpTBY7wMAsjD
lmYRT8nrEK8dl7BFdF1YkdOCg9+f/plC5Js3FHKPekUwiiXFqvmdcXDs0JO9Cp6IR+hXEerRIiKi
dnmh38C0RhyoyJY8/Da6fSh6krVW0TqYcNyTu6vLRukT8TKZ13ofe9x6d3jwAAJPRZ6fQ/E9ntNf
TwZTej0oE4iujfrdvy4Pm7dbqch30hijDC98/H7B478QQxvlEVayF3DK5rW+zSEqK4FuDzNrPfqV
mdKzrLBxU54rAgPxYoE9lXCZ2VFeOTbtbEW+TNRNzWpAKlD1xVX6N4Rc0v6blWFRJmObTrwU6pi1
jxM/UAFDNwm+RPH+b6J3ARzU+hQ3j8HwPBJlJs9yuk+Q58lcyuAF4UJTu1qM1M+myEkiSAfzuHer
6c1RvD1Ns7QTfgY3P7VoI5iDG7T1vOPTszP1o2v/alxZsi/cTlnpQuxj+a7PGTC+o49eN6pSf75v
cjrC2dNlMujLO7l9ad3fwrqCh1KGzsnL5CYOCY2Mnn0lAD7Yc4uAJCeHZvzIPwXOvh9h9nFgnMXD
Ni5gTSne3DvVW1ikO+ElKyOMyyn0cloEa7f5uxetmVjKZsiH9FSbVtl2qyPCM8KH2DtfY4JIEElJ
Kp5GTwX3jPWH+8h7ObGEGIlxrkcIiMl3P7nxwjyIrz+CGtS12CCXl3xazQkWc4sBP5CmQ94p6K/h
AHdcG4nlbWG0eoy0EaQZisrlZBz1jrgLKoN3AJ8MHCIJijWUJw8DrUcWBKFWk3jKCr4CNcBfdDDX
z9KZMvOzs69hs1unQvz5rICVLrOyaonrQ2O+a52aJZ5/kJWtEXCT5l8cbXiVwF+28UbItI6VrjaX
JtazZAXKPkd+fuJ0iLOrDVjqzaYtIRLnRer9QZvK5k/jRjDtUAGyNEfRyIOY0d7TwH4aTYMjQK3O
D0iT4/c+FJg3l3at1h9Eu1Vl1kkdMx75EylC5Pkbc3Sd/espPVOHofmCjDPogGXv0lT2rpYYMF8O
W9cyBcwKgYi01TKrr6NFCJ05IEBGy0a8kZaoMb/8QX2LQIFnTvBHjbR74ydVQJxzWCUtkBWOYU3t
gmdKheLXLTEgkxYRjtR2yUKrM2fTeGa4/ftJOZkRuwN0rAyc6UOmh1k2m30EGEIx3XBTcXhFOeqt
Xe2UlpBBy/wIir9UPtBji/jPKbfVMfSg6zrGysHlSJC9Dcj2X5/UnZlB1FaNYpfXoDRin6E6fiEL
Nc00h+RrWv98ewSFv4gWz0SUnmV/ckzhI4mdj80BJWI11QSHXI9gvSuZEJIXhdUWszpwUZnyPxrK
sHOc31S6Z/pE8SigZVxIgdHg8QC9mZE/ArT1g74PeSn+X2Yr3d0hWpwM7Ut7HS8+wD8IxWRAt7q+
G9voA6x3hgm9YJ9IazygVV8gj0BVOfbSk9lbvkbQ154VVF3vTPPSkS8D/Qn/+fvWh5m1af9E1QVO
fgsJHoF9w1iGzwmMYSkVeGZCz0cRDHV9Dlh+BeyaZF6ofrnj38kzaXatzyLVecrBa3DBc6OZ//fP
KEepsuA6MgiUBfUEcL2SNMEXzDGiAll+WmrBCbnESzzXJoWwLaLbiYmhXVlyMoygJXCNV85mF54W
kBIGNcL3nV7k3r8CLz1qRZRpgmhzj8UyncEnsDM6uPKcXZwddTJDakfAOheCVISDLD/4P8CueBpu
6qXt65BxCIYB9Nx7qOBfcMvC73sCa8NR6jrfs/Eq38mnfSlK4zIPBk8LZj929r+Dl36KYA3x0sPd
6PyDBTktVdqWrtTBhdwCjKu9lrtqJVecoAif/1uyjZXbhkYX3wsdm+kSX5I4kLLx3UKNjeMfJGkZ
IjUWq9UY9orqluBlgIRgvZFXGwVIMhlBh0j5Ql8i2lUfZS2jQtmhiCrj7qSepbAM08UvG2Q/vX2w
iK39ifhHAVNp2cOpNzZ8rKbN5nijXlCt7DR7FUGUJUamqm5NHLG9472S6KlSE2x6Ke54oQm+3Oi0
T3Zok0yWQiOCinNcZDsvRkPYpdyyOp4aBfKqCrPwJCVZpGalmPO21k7Gn8o0E3UOXG39lB1vC9HQ
8et1OX+p6b+cY0Tk7JVsZ3OJK8JLjz7znL2OyMdxK8O8nAOozBaX9q1dUK2iUJDfBwsjEy6+9RpB
cAAsezjRcRq1ml7xqNG0lxzDxK4NKhyL/RYdD1Ddb5ug4qXyuEMfRJVyEQv5RX0VVB2RnGSq9bW9
YQB/ka5TIrwjepBsT02kVsOCFNewiiapeKxyLbcA67jarujxoHemhOyz4Al4NahoU5PDUnhtJINx
Lwio2I1PDjladAln9/COciWlBYKB7E8GI6soWAzPgYmJAEZBrekhYMgqHkTsbZDI+OWJC0J69+o3
lv1nSS0Sap/FOE1nPWUgytkdVJiYm/V2QSJBAujaI9wowUFlEusgTvRCa9MZwjB0APsbcZhZ9giS
/yU4jhj4/1vjyVfYO9AwEBevV4p1tS36sm1bExpEXU1yCyt7+nzie68C9vgCiJAVxnR3GDUJosL7
b3henEhsbAhj5OctmrLKSvdYMhk5NDDM9mVxvknLdaw8K8GYQ8MCNXHei0yg5zUYayUB+JI3t9MV
DTXBkOVaFmCFQ63oxASibiR11zhU/9yPX6YYaqAfdcvBG1TAUNhvCuay9CEWyqdG9Ep+SHfLrOwj
/P+jYDyollM4TB3eCLVVD3Tb0CADiMxNZaxfFGp1pSLlW71r7bxU6D12uloRPSM9UyQ9Bleg2t8O
GAe1uSPac0f1LpQcq+Obumsz8jxRCJR+6Jn8bKXqew10umR6xMejQQPI2h+EnlQSBjS/Otc8L0WG
Q/zlDlqmqSF93Jed2ZjDmEj29vIjLCzPzUMN+Si4TJLUxdrWocWMvnyox5aGyu3FJ+zaMEClhBF5
5Lgqi7mYv0yPe4hFdocWYH+4rxrMLde/PNFvw+gVgF2E9IO47milvLWdpppq6Z9fB7SNOayl9uH9
0NnBI++738HfFIwA+isrzvZgUJjX9FNEhhAY5I3Txnos8jiUrAoFNOLlqdrFTQ6UiDiQjXq/GGKm
FDMjZCMd6WravLDzVTuZok6JEX3I3qnbpEzZapyUzg0KeZWV1UV2DVm+lPz85/wupHI53WToJABy
CqimurzC+3Vsoov+epyiAb0o8wQUV6ZBUXLbjeDxiAY9GMI9WD1adXoGLXnNytowgkZdManlTEum
5SsId1kAWCvjNF3MbshY5TMMxUkw5o0xJiKx4SK/1Bib5WfUNEi8I5MfzScfU0OIPOWSUpsbbIIe
Oit8Ub9znMtckz6f1p2peDxqo+3ViycfMa2iirGh4lIU4LbU593u5YehwACGo4+FS5YAlQya29qv
1ZJ+olkT6zIRVJL2ln2HeDYVsSa7qR0wiyMdRoGKKmQfYe2wUOcQKydzEfQFpyTfuseS4k7Npor2
zgjT3/d59H0PcR2jtlRxAzBeMzIhAL0F12LpZ8/4rRkvDz4VuNMa4n8ZkfvcRqZ26MeO7EzCLCdZ
IIREOgn3p08pEJ+0SSuW6dBu/mOPD5wW4DVvsZ1CMtE0IBN1gGStRkIEkZs9tePwgGJ4dXs/Ui07
RIWBHmgPGZYdWIJYsrjY2nbK4Ydnib3lvGQ9jH/SIfq4Zx+p8+WheL4RIcnF2wrqDs7O0MBKTQQc
WvwIsXayJEStatQEPiPpUaUfqln3GORS2PhOc6kFv3ixtP6B6uW4tgWo3XXuGsk/8OYAvtu6ZWhG
eSFnKXfZkioRsGGbjuTJT2yjhQOklyMLH1ogQXEHc2CeO+6m/FbggNwMILwCVOVC1/TaTCsCATrV
IgL3efANtbcoF5XJNIQeglxqIdhu4rFSrMnaqoas0xoYs13TbukcyY7IjJT75D65jjEalYnEQ7yo
EpX4k/DdhoUkDcfcOicQq+uMq1r0Nt9UEk18VeTSsXnObBWTxbk3GcRG7+v+MzUuExztjpzLYD78
/9u46susB52681eE8ajaFJkmwMHDGRvJgioCvKZbU+VlefBKjUd9lrf3Gq7Bj8K7FlD3QrfAe6gf
G2+9502x7Y2qal6cC3HjBoe4jw2oTWdz5s+tnWGVXBmSKf2jat7MuUekD6+8E36PtWFjPKinpEBv
Pk1pTJSHsr+9U0T9Lr3ILHjDvN9XELu9qnhi4/jdaOeeuzpi2ZcZja0RR9GrDNyARI5X174wDaQL
h/vBckUZ/C++6fYmuvgW59t6UmopK453WvEu0dnDYW2r0f7FjWplW3YLSMVrhArnfjaZuxBSNx5e
hcOeBbVVrf5JgQVWRaBdVKerEYlUC3zbS9b8a+OHGHKhFxwfdH70hUtVVT/kJp8PL84RPzu9zmdI
SxD0jcZ0kbLcLYhiqpKABnpaVkSFRWYt24ip3BrM9FqMtI3Siv5RmoeYk/0lM+V7yPqFGIUrgh5d
2ep5qXCMg8RQWK9HGRNkXEnkjeKeOcBc3PXsYfzP4c9sC0btLL+WLEs3d/bGyFTgARG3mLrSjL27
EVZhX3kf55W8KwKM+R/ttzj/3ZuNRIh6NV+hjAlH8HNr2oWvBbIQGIkqzoQa1g1+W3fOrKZj3S9U
3q8NFMV6NNhLOyG1288ItoF+XGrvFO/MyeLkpXg7kW6NbcZKTMo0vwQ2QIYTD999dEsWojYnWIEX
TyzSbyUtTk+LbDlUtsIE3NnGCKzcR3k64PtFDrfLlxoo5kyovZc35rwMS9YTAakexHQpMrACzeis
5vdYqp4Qx9IJSH4jiELflaiDtwapjBx1vjclbSGe7VVfmBnpgcNUnfgjo2PHSKKwbOu5rhLBHKgJ
xyhFtCvRGRbooYpDtp17PW0RFQod4ao4MsmEvNS8y3ISDS7Uvze5+IQJVXf4oep1wGtSOFWZSbcW
mn06pQH4olx+ll4CaZ/PTd5came1/mbkWENgO6T3ySqHfL82+J8jqxAizwRrKe056vUPezKvNhuA
KLJhAmOB9rXoFnZSTZzzcEriMFhgzGA9cLmGG6RveOHFwRoDhelAfv1WEnVFySyXSQMMYZLdzTXZ
+Zv+8ge7wkQR7rDRos1XsSQj7YLTewjIdECBmtwsinIR+/1t16wcloxYvWEvxO98oDo1jaJiUZ4Z
zoQMgUt5JydqliR5RarHEGihFAPUUATgj/H9vz5mXnfJQEidOE0qv2NUC2Ta/liQTZs7ldMda6d7
2bTCVQ/Zodrwlnkhi0KinrqdYRrq5Vm1e+Wv7/2KFkIyzbr+WZOwoaPXizfV0ACQzyTdOgDys+KX
SHVurDXGTDySnkd6dHOlpjXUMDO4faQ9f3ZBE/y7Q3aI103ndFZY9kqJvwnEY6I3DHtbfEoABqPE
qoGW0SHWcrWJHgOvpKts3+pPRRJz2ArlP3CCt5b0U+fw2FW2ALNqcGUO3s3YhLFRX/9yzZ68WSXK
9ZWkOch0btQiGaQgRwzXyVvYy8NxFTKXXMGzezqxR8MTaRJoleWfreWK8QbQqanv33kuXGQf84ST
Urjrr+UwW0fv4uf7oS4TkgtDkCYeZjGRJXOPZqIGaEDaQBDzIA7ONhG9pBzD62lG89zNrrMKYZFc
F6XCFeZj50smst1gDuwhL4MUgNO5FTwPzY6x2tbDP9uXOCbL0PZ452TN8GGpoaHGiKHNTADpZHNr
SII1o90HykZRiGhYESHKn7lwECbo3UeHQV+j1OsKVeLkwlrBChFH+4dlf5dLi+5hNSq+ajkD5/BQ
/bKwDYoysWci4JhG4iUGX3+FCUr4lkwJdfBo0zHoZRH9dNgifVYUozNZHAnM7o2CJ50HN8iiIP4P
jL6OqNxxAaplUC93DkIILMmb3nj/H7S/BYyMwtXp7fUA2uA3XRS8k3egGDnJYnwxW6Rx0L1Sd3C8
hepk3bMMzaWCz40BLp+eZ7h2Ckmht3g7oz6xOuOl0mX7u+p6UY6hRbN6XqVPzHhMXoFp0C6lEz7p
Y2n6Ugj5VH50Foq2YQYyx8XVbvyIRNXa3eggY38NqE9JFDhBk+vWdAGZr1T09TdHAtwqbIoYPGh0
zRbiaHRfE4GsDvWW2HhxDAA+Br7pCFHcMfL4cuZkV1mjXGiaJI7vn8dDFFyobsnoVS4wEbu3QlbY
qDARL/Njyciq/mieqQB7EVMjCpdhXcg6WsnNY+7RlpNboTri4ymHRSf+eQpecKa/TH0qTIuGbQsi
vKJEoznrBd1483On1krPUGhwEK1l4gFiMrrSx9k9JvuJTBYWjkr9GJg/MhgepgKk9tK23EozqgBZ
ltVky5Jx/f78+aqoUTCG8u5o9P8SmBpHm2GKYf+JjIQmq6X3uBcJASDOjByKa3uZcm8bq3REDRwe
AUnDrk1yKS+33hkQW6NNQMnwfmGsJwnA2d1oGkc3Dj9AT+BoXo96UClrp4d5qRIdqhfaXBfqK3ii
osX9HcT3ySHrGyVVKxyD5kzPBUcxHgTxngUZcV0xwahFju+MhaMLbd6tmZSV5O+F2cdgDOL+i0kr
mdOb0A/2J5t6m2lUULQYgwUaWKlZI5fzvRMj7PKPq+Rj4ef8z21VnFZiSUCWTWhMkX0ohwlQh+Z4
i4aNbx8UMBW748aps7kwI2YZ8ZBBaGExQqi+Dx6XG5PtaYWuAa0cYA1hcCXY3hE5xSW1urtO3fhA
Q3ECTawrI+gWolA98q6dX9pcJpqO0ubCyQGwothnAZmrunQqYqJocSckWW18lFYTTp2PL9GhSZyh
roktMwhT1y/9HTIbAqEYYhmTMDiFBsC4Kd62VYjbcLbRequi06BnKkVxskjCrqxMfQgEPd0zw+oZ
97iswL3YwDmcF4ic8xqU4lqY5QtW3chvRI+2KTxlBS/r6+conw/cXnHuEK90+Luea9+Hy3SPn62w
zWHyxWNo8mKWZCWXuV+nZL/kvvWw1rINPF4YJeACAsP5X1HzwE05UiDGeeys1talw+Ievga5u4dL
uHGQZYjjoIJ4lMtTNn3bFb92FbSxn0i9y9CzrbczKwb46YCIqbka0OOoUVBe4vSG4a15i5ghP1nR
EZjGnYEMUt8oflXZIntYMIygKc72cjH8PoG9lVXySoMPhjaDUxxVZrR2pBvmz6ize5FSCtQJePF4
bsyFJKJ8AS7Y7oZSIxzSKMfXrbUUY6iYnI0iikc0jX21+HIoWoK5+v2jI6+dM/HgWh0DJ0fgWtt0
WBhIl5rey4Mh8ge0gg3k7A9aTym6/FxMCoy//+w7oIY85T/lWrBbWZmtSOoCAQYoY7UO5aSrom2i
Fnp3ZuSx/D7h12/EG1qQA/7TLKZ/fj3af1oSneJ9vitrDk9Ne2sKLZq66IUvBEIbnLmN1T2ww20c
bRKqP2LO2SiHvXZJHld4S178CjmbMv8mt265bAiAGgoKFgf6rk7Hp7DgVA7AX6PgM7RY4EoYlQFO
gztbWCIA5tWYj25qnw66BYOIixiJ/LHN+RHYieINNjLLJVHzJOzxZWYqIHGp6toEY9hbZrmm8m9t
bMHWQMH1HrLZTcYev2tZAuTZeOtBGdvp+RklN3vIPM4hMAW/0dgtl8rJSlNG0V7zGEEmbtT/GE9y
Zfh2RYWvIg96VyzukgFbIJPbqcKetQOqZnbSYnAUzKAeV4xEI+Sud4fKm2ZbTwrzfN5ozEyUjeXt
VBvO8jiNtfjdPArxIZHpeTizTE0IUNgge97mj6h07WGyxBuapgU2TXsAzLAAr43h05sY4bq/rOht
aHi4VK/6nzdR8PByqY132AwO6xAgbVgSy0JsnQll6xacv2GgW3jra/4GFJZ6e31B+B++1pZ/Rxwm
XK2hSVHLGJpwif+fm+5S4tmfS3pJOzN1bjtKfHkxDbX0n+r+vyfD5wbQTzXZL3dwm3Da142NUVcQ
SptALM907VRHToBhKc+DM2PViDgPgWxB+APJay+i+fWWg382FnEVGt4L2ouq7VxDyVkFDahj4AtS
uI78w1ZKGs7NxJVPnUy8CK+Q3gKiU5AXhulNzX4W4A+iHZ2BDtNWYU7QVogRubKcJidYXXR0mdJV
umicxYxWhd2MBuFMP2lrOesw4FSL/3MEVMAU2t9UiS3qwNQc8D40RaNrd+RTB5OE6X7k6NMOYkow
ugAgTBpf6V1CeQnO+83I1QgYJ6aJjNaKajUPY2VeYzwKs+YvvNynnU8BQsQutViiKnh/ftoE9j/8
9/wU14BI5bjyr+JLMlHLrXkQuFrK5sDSg94kTbfOnBckA2wpYIYjwZY2kqrwQBecYWbYRZ7wuEoe
JVyV4EqYaIwEMN2tj1jNpdBPH89h3gOOduJUV7Xa4Vhbc69W+DPz7DaeQH5nCLMrf7mIiQ7XglxU
wo5iev9BoQeB/V16lw6OdVU+AILLA9rs1/lju2v7N0HEiRg+MIntYva8GzBMsQ7rB5Kcr/INTS+j
R1KZ8PMXq+mgN2TpKQ92uQDVFkXc2xWFw9/jmZps4fwXzaON1XolaKm1o5LIo0PoNq3vOnw8FK4q
TsINybuDJXXP2zMxu7wDApr2pNVT0sOPce15q44M+ys7g+h3c1jaEgkfBvvD6PyyERsWdegxnJc5
RMmsI82q4AXr21bvFGF1baxh1DivEgy4qjuNDbwryp1P7ZWhbTj0TIVB0jDiCYU7mfhpEzEo8is5
/1tuSZx3QvLlT8Y433sVOjQ7IcolcQR/cKT/sDpj9fJ+qsMYYAVKOBd/RbuGNz96uyyN9ZKnFchZ
fyzYNE5aLArpZ7XF5ef84z/ohSB9GFtekmGMf1r6j/9Z1mCoc9JGhkpaf5yU6JBdkapcgkZ2NRRl
74fdL8HcoSlUnIUWP5i4VzmUjABbs9MZXKrXx5rH6GwvhPB43sp1ZcX98Mr16YxJqTKBSb3N8oI8
BfSLPDHZlX2Q8CvhvzP6e+eVjgINMkRUfYFyWVq1ASFGWmz2bKZg/8fytQWnyDw0fDVuiUYVqjSP
sGncg6yEV2lYIL6t7hrB3Q32pwh4XzKA11EgIqYqlHy/J7aJYMFKLokJEIz1M6afoe6lrpsHhdlE
/HV/1S/rtI9pC6mIWm3GA2J1T12jDeL02fHJMbZU2xoCLpBq/o4zmAz06YrnR/TWOSDxtaKvzmyp
IdRRgbtoW1dzGjBbUEmRQd1bC7qaomWXZKwCvAFt3mmd2+lxTSxbA+J9nFFRhi70N58nRBqaoVZm
cyc8gMLhiAe/7BsmIoHILw1b8J2Mc2+ie9MVwf3NVoJ+tUO6zu46pJVHqdDLBVfmuirLNN9iP9rt
cxOcNq/U1dMzx8TzfNy0lFDc8zZj5b5FSeWyA27t5hlbzMo2TyE6Pkd/gklxakFJOs0TuZVEQ8Hn
exRueEl6XzUOFu/eKG2Iq99Z41HYf9bZXUTShVi7hUWLm7H+/l8yanvoLO3KuiH5YWr9pZuVfYnn
d3QnU00eQCtcBlT2EqmKYk9lDYUD5fGMsF52vxC40wR/JV0mon6T8L+SFmYeO24mvDQa/BuGurxx
6XzbnmfYJzzctvV0OK1cUJya/6kDGXJ7W85/HdG1asqlwTUHI0rO/6aVd272sE1Md2PQpnJTwbRf
c+5yutmEL2Ko65+8yCV4BoyesN3ox1qX57Llxh3whgEVCt6nIJOMJ+sC9yl/OlOE3yepcnXpDrmt
S4jtM1lLJsj79Dqp0l7+/NnskdSF8/9FJlNB1V6nZaD8iCQlJ6S28If5D/6cMKBfjQVdpXTQCfKn
gBFVM7d5PX73E6Ske7I7crw9Y5XWKLtcjeDNiy6WBjzaf2KTEHBWN+hTFCs6RESyx2Xk1JdEHynA
Kl3hyS0jPy4xii6py9PUZTnlGYU/FMVgHbiP9LBmcD471X3d4iz84O6i2bNwonaSSCmvVYusaVtd
Jntx2LP/MInoo93EQKwsuAFFHyF1YAA7AIRESvad0TjDZAj9yXTY0soFfwH+D++tbDkMZNv1UX+W
pLIgQdQC5DYxNpwLu1bLG68oJC3tvvazN8xCF1/GCWjbemyZaxqamvK9c1OlApbGLUDdtUIj0paF
GnGHmTCAmJ7FZfbeyNp8d6QmonfUAQhVWBQ/n7Qw4/T/hstpUf59Qp1WmyjKajp6gKypydIKAhnb
3d2/A7UR/e21zcov87s0Wh652yRa5UA8mfriUHBqfNRmA5/9NG4W1OzTkbC3XlOef5ONzBSnXDhT
cb32n3c7OWMVusnR9en41wcnWbXtxjNdg5xeC5AlZv7J6GKkweMNuQlhMvcGn1PLfiLvZ+QdpaeU
rKfEdAaJzb8IhjIfBlUuMRD04QSYuFI2jyMdEMNmslonoREvHXDn4bkD0OkTYe42ycFSzwHqMRMf
NjbRrxI7cl9riLdgbngTrJpG16HePZDp541/HLtztuXhhVa2BxdC+00MSTzLvXJlOsJg2kqFoasx
K7EsG5ws31Ri/lPvvxUTlpkht4KC0CxV2CF5QBX4vLifoerKD2Go36m0/nycluy/Ff1K6XGdhFMR
7c0n5c4H5XI8rB1P8p1A9CY4SnRM5fQ7q3/wSHQOXRV+4zlJtbls2KCiPSnxIUayl243ssYnzxnu
uEsL3HGYxpTACNIurInVO7hKG8OM/4SKADfPK4h3azC6xmmywD8MAPy8xx62xSEeiC3xKje8B8TC
sGGghd4i1FmMEAZciov1K3+LSAmFHoRidcTHwR1jFMLP/hhM2i7+bzOxi7+f2R1VfQQxlO8kXj9+
F8akprJHINcpZ0nCbibAaK91u5DXndG0kIAfCahcw6HvLw54dn+ISzyJAPG4WswNIgS0qH60oRP4
cPnV1pYHayzrhaKmfhWTmLD2Wmq4LwfIK1Aomt1zqqKT5OMhlN3hDfCpZq08p0p5VM8w80mTJe4J
ZrgBeFKbZsX+4r8qMgMw1kS7fJNpxO+siec/wGLSzL1y+OAYjbwII6S7IDqocDLBmm8EBZHY7nun
hrCF08kgtHV38JVCJn7Vgl/A+rkB4hQXJNqvYsz0FstVQ1FeHJHTe484VVFJw9Hgynw/FRJREeqt
iqA78eXGvfKtJexbv03oVdwFY6bOrBs7DciFKk4Xn6FyqlVhi9hUumnX822GvHOG8FQHr0I/vZ1C
D1Yq4s1LyQLp1G0CyL2Rpyzs6WGFOOFOjayOCkQJ2F7AbJqKbFptYSvi/STb96Jam4m8tYkGk0K7
qCkbSW/DG4iVbi+g02zai0QLu6DDBweCiKduFwU2eMrre5k1fw2eL0EQNCbgDhliQQ8U/4Z0EJ5I
08L1w7Xb1GX53Z22fIlgXSwJqNDgnReyP/oF0UQqsbYBhlackWMqkWlKrkKuHVAlk2W38KHsRXJf
NdhUEag5UppPXNlALeWBxp+lyvvkz6o6petg0LUJw1ZB19fvvbg4ut3VGX8pUQ9psLzYW58dzMif
R9GHPfLR0Sxw1LR3B5usR/KhIo5ECBbEvY1CYxfIhEcGhcnI4P2FkJISsp2voZrNN5Ad2AMjB0KO
PDLzzVxYCgnskZXoKvN7w89qQUPzW69R8iYibeg1066lbkNlytDXy92gjrT7zdDyAmLKRN5KPB+Q
MftdaXYfMy7AVYujfYXkcUvbt9UJUqfISWyUnMdWz12OoPmogbHeG6NVOuuI/l7oNVfBtw9xTW+e
yBFQyCtTijIHoKhG9bcNZieOVxqG2iVvPfEzTVkj5YfoFx7C0Kht3dxyQRwXYescsTdrB7zVqIqX
zcHp1mNyhRdY1idhIVUmLL5TPj9ldmeY7iZnENL6no3TX5tjbfF8I/IuyEOZaziJPW3HfMrVxyEZ
JnnJtqsu9HN6XotSweHcfxSyvbvnvnpNz8Xe+Vhh4yCDB62pqpwnX/N5jO0xhy6sp1RvwTYAVexd
PmMLintmS6oMJeYlAqria138qdC9VCIGxwsBbjZE7nryOKUBbAVEd/OzNY9LbOnqGbMP6HK0rq8s
eQ8hLCwnX7K1BvSOJwBm1BMlPkUEuYR2ad1JohkVUVt3qkxQiyu6S/1QcTxtKWUoe/nkS6gUTVz7
vlnZrsdCebNVIagfcJ1S5Q5JBN4Or+u5yIMniqQgRINEaTYqCWHzt4Qh5gcPVjIn8tnM6hpMcU+A
/yYH6Lad7tOrWqQtzNihpzCP8eyzb/j1OgBd32cYtgQMW/CQRkT/YCUM5gc5jgM5jfpi/qN7qkbn
q6ox5FXytdY9eUTUFCxAEOYn6kbD0IXrp7RleD9r1PkjLVg8L0QNp6sxmauoGt7OwLMxiTZEi/Ng
IfXS52QHY6MDp9SMDXhCJsC25/PUvMJVN6+loU0QS7GWeJ1+s6FKdgas6HF3yWMH/xwyuWhrqyC1
TX4KFvof1LtavM5rREkaL0ejxqBYmRHUSpxLqMT2DFuo6KKrpzQNhiLFaKXgo5EigASSosBx0ry/
Xcy/8Vohp3gJZ8KQRdh/+v+aRhpse9NNObnn4loanuGzsxsaZc0W8gCB2r1dyZ7zmvoEMOY7vXCz
+CSeW+xTIGyRbDi6QU8hJX0Tc4IIbmTKBS+OhUHmifYwS2Xq85+JQqBeZ6tgjh8wxsJalRY5T9xT
nT51LejxcLEDk4P554Zv4OIR6t0Z8C2Nyp7JeNbLoA8z8ylQ3uih5Da93tIU8c0uDS33Ze/nh5qH
+06IFSaUs1jA/cwCc/pi05hcBAFv02hCqRQ/edt0Bi1HPT/fXwcawzo4kOUyS4bmRPjbGWlymEyU
WgebRrQjl9RLTmUpqEJcaHehKjpueFX30I6+kqvCkxVVfjqNpW05e/Rg0q8ZdMdEIr4wLKEWPgGt
gkKZDl7wedk4bPjYQHFwjlXDURr2VN4igUXCfDJCcPvyvo0ZjbM10qYd1HV4feWkCLNDPHrUgrSv
y99d57sf8kWxIHj7LIP9S7Di4Jzxy4su6S9snNk1wCg25iaUZGTNGFboII/JFVu0Zy3i4/KeStMD
SKbYfEWBOYvoKW7UAcobm1FDQu5nJyAQbr9CxOUK6bfzSvGt1zxCuy5HbvDqpejKIUBLui2qhE16
1sCY/93PP9HkrRb/+JZ/ZGxHaDMHBOVXd1C39ilN+hX8UQE0G40Q5GyXSRs+oaNqubKAZ+uSUaRG
f+BvhMnl67UvPxFFupytZ4ro/SERduyLBUDY79zJdVNKmVNZQ41jXipMJnq/TDHBvyON6Z+Z3eUG
s+Xdh5QvmacVLTK1BOcyRQO+3MfBhhGBbC8c/+K2iBPSvJTjJ6GDfrOtBb23O0RlE9BoKHbKSR/E
gW+gCu/xXTp46O5Lj/3WKqh+QS2Phbsxpps2ospyjZMf2zyusDWohggXrjbAwmsOo4LQrDDl4UqH
DJeZuPfFl02sy97psxdpxL9JXXOmbICvqQ3/ao0LdW5J4Nu46LFPuotQ+tHQ+2OR1lf2uwTbAoY+
ENGYdDfRrNHxVLO35HC2hKbyARWMwMGAe3BhLZJ5W1Ozg08hKv+sA8ToTsESGB6T1sYZwKOGphta
5U+hjRzM9NxTZ4BoMpFmcM03+LfoWomBa2bNpSrlxhLPzorGZmNEstgQ8DNaAheRz0TrsmU/WEGI
7Eizu7mj8Z2zzKlqtg19+tYzeAt6XAzk3FVnN/5yA63Z31fr+wVOQdRYjUdgGHevmu5SvAXhBl4T
sb1DWLhmxigKwzjJLz1MHq/tWXtRVIku/fk9wdLpGGnx88nXIl0uzXC2KqkFtnPl+M69f7wpHqVs
oet1dDuCr9jERT/vMNQi0l+tbuFSfEpyKQ1jsUO30lSJohOqgB4FpiWcsKUB/KgIN0PcXF/Ymzou
0l0NXonJ+QhmjmGubuQOLDRdlLB4fiCWbOBGBH8DBbJ7VrzhbsR7aHyyKw98Y9DGqA4sW0w3XwWa
ff9Zjl6ey/hj4JHZSuNcac4jHHIttOLtiON9s5DHTxtylNd+yumJbRVK0F22m8LiL/ubbwzLpoD2
RCcSJU5Xb0IoFhFcwq26w+nEgYlCd74PcWMs0qXi0eV/jdPI7WyEfwLAdmiAikkUU1EbsEvmPbd1
njJlHgh9pgCqlGPl3rDkVsVmWzpUHd23TP4w2sOIvkuQnua5Gne+S67BWjEiejn7+JXIRjqgNpdg
P+AazaUl59PPoRTu3WrVe1kvNkgFxIyNRi7T53VvcWSfT2HXKXybRwFXA38oSwNhff2RRqcObLLZ
N/K8aMiSuWTaJ7Cm6U+lmeEogUSnnUbL5TzCquNOZwAEhj8CA9K0eMg3bHIhR65i/fFvKfypO5na
iiijMbo+cTfLylnm6Q3oymBD6kK3fefz2GyWcY+uzXHv/pif5Nlpd+BUmzRNK/yk8pwGYgW8OYUc
BjpLbgYXZxd7gu7gSr8URAUW/1KNcb/nLIELc763sZ8UwLC10FjlVEXsSAuWMwYvPFp7YNzXd392
Q4YBk38zHLyz0z9AZ0td1iYd0UJQLohI36xpUR3m1PeGN6mJtMcH4lvD8L+/MymVzny40bkOF6zs
YnHHE8njSQdGAoIAnGqX2uxsw9aZG6dpb6C2VyGA3aiGpwLgEZjWs3naSxmewwM9/rBa31Dam5vV
LjEdvUM8Sfk68Rd4JfTjQD89UhTDYgmCjY8W2lZ1l2gVxDuizzto1WrSqlSHvV60SRNITFQ6uA8v
KZ3fM208aYXCgBEhk7fTbNx8R8LXuC28ZIagtPz/i1I328np4WiECD+IDcaKPkM9dWaBxP4P4oBw
HLRU2VJjDisl1msfiJdBbC0Nobbqr9Y6FMAN5RFkN4KnhBdzvfeOMTkbi9IBif6AJ3KaU+R9lXBv
POe7AZMgS5Mbx2Bl3EvhCFJ53PDoKeZ4dusu52gxTw1i0jfWWdLYTg+e6q9+K5Uf64+bpfAfAE4f
QNTfepw8C5ViZg/9uWksH443KyaaimHV6TuHMSzVIQNycrEWnkXhfS6Yyyi9wytX7RbpSjZHUDti
WC76c7Au+ZnsjaJVvxTJ0ll4DKiMc/HiEkNdyWqb6tY3qxsVz4XrDqEb1rudxD4yJCl0fAwJV4tV
MfjhZ1BcNyJ74XSFoarWpfQRqHWBypQN63g1djkSKzfo/2dQw8zEwY3ttC/RAfLXQIqr0VfXdre6
zMtPRsx+myQkNx6DS3aUGq+9AWv2lEMyN/WKIls1jNjAYgqm2+0DNt1nHH3I9kQwqwqK0ZSWCrNx
COgn8268Yj/NPlegxvbKxt+YJSUwPQraTop2qJVZAiXWvMwMPTcJxbtCmTvKo8OymIt6asFzqI16
2NZiNXK1UnZ3K2uM4junyKnfTGLqtAu9t7oO9aaNJeOdwMgsYGKnoVEnhsKaG3YG5S1zANk+NOQ0
Cd4280QqtLK5+V2uruEkA1gi4yEqDk3xhKNxVB0BlmIYbKsM4xnj2qelIVPBhTPKP7VwbWDeJh8c
CsxKlCa4sKqP+NG5agONlDClTSMAS1qDCA6KqXfTW2bnuiXHm+alX4Whfz1hbh3LlZdqHduziw4x
6fQ5oA5w1uFSxISTUKISWUsmUT2l/MEAVzzwpvc+9daFp1xE1fOGRVaBLP/FKH2QaEf1pCli3ZJH
99LtIC4hH60kPVMsjB7LJbkaDgX7SLmQ7bN1tTqBR587guLVDFJa7GAtVeg5vzUEx6IoNFZAgqdY
6sgmuO0NyDXYWR8QI+5FJk7CX7fCD+U98VjHNtRVMBU82CULmkmYggDaU7k34jXZfcw3ZDCnGKri
Bg1zXpnGTjNvV2U2PNvaXu3WYqQyag5zDT5Jl+iiLt7TvUbYZPlWEiwowf1TpNPsPRTK5AVW/PcW
ZgXoUYSymfOfakJJUwHICCL4YNN7kd5UFmbxEKq8V/NyQGgKRw533YV/o03GNCiAZ+0PQ8aRl5pE
q9DwpwU/L4UehfCP/H9URQKlqeYhw+fBo+ZOwC62i5LJVXjIpmxEt4vAsSVGEBNdweBEpZgKxjcH
HRZ4OB/DvggeuryUGnsY/9CNSbG3L5O2l4tanvbQs6WVIGfh+KQFFNtyfNIDuGLV//cuIrur8EoJ
zhjaIdpf2MfpL9ZTiciv5HzqZX5xJSW/LB5gUWS3rE/U6KRaWvmPbM1EiE4h9WTZPxNk61FUNXyZ
TM0Gu4JHbLtFGcfcTGq9eQJ/jKhQG1OAMtokjwUYYNG9icLekxxmYVZnKNxb8DQhQVbMvlXmnBAo
X6ZJyjH3FPmd1TjJv34n1q/V6gEGeLkG1DbzZBfmKdPtAt0ArhXJMWMMp9h+QAsutu1aDTTGCHcW
Hs20sH24McHE/Az1g/b/fR6+bGTE7OZ/C0kZPVRG0Xi3SBF7yPwr0BI3xGT6yLncBG1LOSlcGp1j
emtSfRMxvjGXYCOBEgz42MIeA9pR87rlPPIk1UTajkoa48kVaO2PfIMo1LwD/6P0tRL+iCnv7+MQ
bhTDBfvUbRzCMaK/fGC6Z0ru59Gf7JTMo20dc7D7cYTnwmz0oIjhR1qOCRG6K9Uha5fvtLVVXxRc
drrDqsXZ9dfnPTVIeVadh3V1goSn99XnXkFNCGe4JCdXC9grOneBGOeEQtzoTfjgYcmXQmmYcf11
lgm4BDgaL+cpUdch+RcvzPkzN+M0HJmZRaPfrG1HZ41lJ1xC18PFdYkLppsZLC7TXXZHINebzA2o
Nms8xHCcYKx8hAgOjfFVkbcZVRrVGCmzEGQmoTqbTOYLlkVXysArhNAFyVQg60+p11AGsZ2wyAk6
jo0jiMslArNHyCrTCj9E1FXR8Tp4WenRPaYT5p6tnKmmfgXHkhEBd59bW1TSTwJQAss0jgeKDFf2
lm4//MhTRGd7fmgqmYY+KWEi1oRT2Ew25GgIVlzAsLkGHuqDzuMTxfl0GVYl6JOAPZFkWQvERlLL
Z8crsSyHWHFSCKFnVER8oznDU+VzMWWGs+LAdlRK8B2LKYznYvrTgGeqQ0dOCMTcrxA2AxRBp1xD
T4cr0LN4MRKFKrAE2dA4mZdVbwONWP6Nsqlh86wNqNVeX39fcnQam1oUI+BTzMvMcoANQB5/svq0
VVtjPsnH/tUk2G/XPjlNN4CDvPqGaz663n4Ems6nzcAc9jUeTUD6kluAtyFUC0iDGnqBVfixGEYn
a6SmZ/o+4RQyrjkpb6oG/J3diSK7bN1hWSFcVIbQdS7bc9zweM1zf0p2ZqUpvLMoOPaKdscagWN8
5cwct8RPp8ovxncDCGiuWdzxlRQoCqfy8F+MoSh8sFaLk3/nsRtDqUgijrtoorJIAmIOLEpddfqa
y/XB0anACpL2ZqaMHwfdofwaQYePo9/1of+Og3FQjLluHXq+lX/XDNij0x8riQ0RoQ2s7RuxZ73f
4konNJCXjzNBntOxt8z6mgPd3d2nxfrFcKbklSSW80nvuwB5OAuRGW2i/sfQiusUFugyCH8JKjHd
6FxW0ZfTe7YO8IDLDPWtd1hs4tTskBgtB6tIV3XIqeCmjN3WPZKKUGTD57pILgFW1AH+4oKAkHps
VQg7OnWC7Iwd0PK1NehdQ/55NH7d3VuJsjwYi5D/zc7qSqRik0cbxm/4LjBmkp/3nyUJrrU10ln/
iccWJ466+em7QvUudVbB/nUf6ntfmWqzeDpWV01crh5iAzhmS7O9en5RJ8SMVA0MzocXpvcsqezm
H36mJ/+5m5v/uYAP1JUNuXJYcKtnuKhVqN5WgYRatYxYaUXBQ1m7NlsAehu9u5ZBlwJLt6BIw/r7
mfGX89Xci+SEptUFCKWgSk4/l3cIfmnbVchi+m0uH13tlqLw0CRiQyl7ayBkeYa8uVpMvKAc74zD
vCv7AvpeYm3rfM8k5+6ly2cadhHG3LhV2Zc7GT3cH2k1oxTt3JWbGv1NUBThzoqAaPEh6rf80X/J
oYFZIRW9V6LDEgQZtYqP5WIzH5acbi7nNLWv9zpQjekAlxlg0afucbrpVMffWq03AlWnmdO0uGdb
6wgW+E+foOQpGWZ+LyGRGb6vZPi7pufbKSpmfNvwmarbWKroJm09Z9UF0o3o9/rkEyg/OJFLeXyf
OjZfJwUVRHQ/9ZFapudM0P0hEJjeI09sKUe1OC3O+1Cw6OiE3HhinYQ7w9Ev16hkzANJbYtT0BtY
z2beNaHiyePu2ulGFWXEhewbgggXN1z5s4HWR7oD5FfvNUj4EMLD4ot9fGqoYxzZvRWBKXTtUENY
DMgjBin0SMDWpR8B8cK02J3r+FwoIG+jLyeWWbCpiw38PVwvis1AaAQNhlTct2IiuMtQ4xgTF8sE
aksoTGI84VpHTHUfgxlYsyfvvxzPNkjh1/YUPsUgR3XRlJOqw80R68LGcAFKEfRJtkF8dgiZ9NSQ
3lCRoQFc2Gd59Kv1a2w/i+cDH7xMoXDl9bcqPa/vSvbMHkZvTy7Y2SJVZcBrumKwi2LLqsMILwwB
QLXdwEtV8ueY3Uq9x8dLnS/6g/fKR40qGEKDMNVm1Cb60uSvyDmgkauvqny4c6hocSTiltTqiPxr
1MrNTvrXHEVn+ZzYUo3os2V/m1rE0afwTuGnBX0FNLaKCYPE2aghCi/pCTkP+RbZeuGYc4Gqqi3T
j6Z64XjTdLO9fsvGFCggJuzeN9GxZnUcVtJNtX4M06regQneR9WEy/0JakbANuUwqLenSbj3LEpD
Qemp4OxwOfnPgv50pmjfYf6BP5QooC5Y3plXIhEEtPK+AJdX580tsXUEQDZwkJL5zLPWzS4EPPqt
RXDlOXk9nL3fdrQqWQa+1wn0AKH33+S/4PGJILNEqjMrxxjztTxGW8GrCwO1L6XEOCyjoKFofcqz
0RWU0KpOnvnvCXAtLyM63HXqYKmoLDts3hpXY7qCCeqHSvZW336Bc0xKsc9JYDorvlNcaaDsDZ6a
xoLxemsteHSF1qZjUV04T5UYwg9i9Lxd7MYrRjXlX9XQQqZDuz883qTPtqjp3FC6dN/garVgA8bj
nmf6XfKki3Bwf0q98dZmk+rFkMFOkjV5R+nG2Irrx6TXbsg1n0w3krjsMODu47pDq70ogMgqv5j+
D6Jtz6OiSy7PIskHJxzhSpIQq50D1V3ugDUs/+WdFOuNwwZJi3R/joN7AvDeB14s3OrWvm4Gxofy
fvvd5OXQ5qGCIvJtnacnoz3QCn6bS+btMEehRj+6euoiY4Wo6dfJamDuN1R73wesSsf6+XviJBhu
5pOz2MecxGF3MrRGiYjayOn1jb+Ld/4rkX8nK5LcFjUdxDCazAYSIUdlR/wG6oF69SPhVRhlajiF
MBND1Gc/v3x7vjEbB+8qLH+9AztN+7L4RiMNkJF8xj1jgCct4YLHXyyl69qiB0CZKgiqz8HVUScn
+R4aw5tIjtjb1qubxBpBQrLY12mz5fyybjnWwSoT7ig54ALNYWB3IHuImyGJcxgq45zg5XJraHmQ
uoCBMl0/kU4Mp4JatBUJNWEmbktfs2dGlz8omJQmlJuQuExmUJaROjf/Dl8OA7P6rjbWkrRJhsDN
iZTV3fcb6gENzAkANWdmE89irJ9dh4p85/wt4lc8hRIYfc84AvjW287DJTNWQdU9k212KvZk/db/
D1KuULZLidgIv61hDFM00ifpYxPoNamrUnfd8d2ziPvdX7qvZkqPUC+vTp2sbZBgp+1CQBgE7WiE
rWhcMWE+hJS/rqcMxOuIT2KMtEczwlBEB+HZGej1JTcr8ZBlVm2B+zNC32wUnLuLt2JTUMXFbeGD
PrwKtDTLA0/sXtLDV/RtmgVGNoSvUjMihGhIClZd6U+oEys+EmexGSQ7OIlULGIV9uZEJI5adI7r
XYXmvMFTHrHNBohG5sxWwcdn6QmGI/mm0vTXlaHEtmRCpnpQK2lrla77y+i/9dcblw15XZfceRzn
/GV1xeNTk5I1/pJL37iA9x6sAaJ50nKtfszjdCmdlqLFwNK5C+321d1A1d4btUoveJc+I23XjxR8
OiO62dgRJx4Z204HYbJcmJHTpxj9gPyavzgZnDN9WjNf/DAdtH2aoyxNOtB60zMzS6y1n051bsUT
/OA8NG/SQop0ZsfDGSrsdzTIP90vkbaIMByyMPKM77samF8Bf9aSANsQ1s809PyYDURacM56r3hw
JmT99DAI2hrWjAJ1VO7fGY0IEPex72Qpkc8SEiO2SCPG4QLPePxW93jApHkd8jQaInfgz4bBEcp9
LveSNDf2OwCTn8VK3lrRtV4iq6H64QKk8a45EY/VdKyJ0YRk0Uu/xeC+WlZyGfdmks8Sp2HC6Pfg
p6B1u4zzAu3IyWWzplVrr++Lar/vkTNhm4BNepdzKR50vlgCrxQKQP/nqvnrUDJz43MEFeMlwYsU
kUv+IsSbhlRHPyncZKgnnfoAgW4HcO+xcJmRDBvpon0nE1M1VzQivdIfTizlcPsM1n4D93Qnf34g
Y18jkwOvvpm4RlIsCCQQXkimYuqCtMEJANVMiyWUL2nRpvGRbVz+mOiYYpkCNeIFpIRqFzI5I3v+
heN6igOeYHlwmwWq85PKIbrPHPclBKRoSo1qpDrAamCFhSy04ZuOi9oZgev9FHgmtnsWl9CebL4i
WZTiHAJSfVYo5AaIN7p0l76sTuz+10gPIPWRnGesI9AYFQfRV1q1ixp78+Vu6mVViXL3oW5fZVyn
57i51EHPitaxnskN0VoymQbwHPWdhlF22cp7w9Byd31GFhYj5Ka109UI3Zvf+KIR71GhJ9f6qkOR
XI/0izHzUOPkezzWxvVapHZTloCH1a8cJKoZWkLQbGQse6xQunnaRLLz9gZDWA9husw0zn1XLIz7
TuwHK6Be0VyZIuQX/2h4J6TPu3jltB+RYk4EgDvXUn64VWJeJ46tol7dvDcrAv+XPb3TjNaWVycj
C9qpdZKkgwXIFfYnprRoz5MYbsp5Uw6mnJDn/Bv8dyyEG4Y/8eG+mLKVxS7LXiyULxmdsZM0m+DG
IU0U77ZfVDT6g96+DbJMp/bCkXSaDLGdomdrdr5j9jUAp9NScai80EzXHKA7jajMkR5lCRoEVPEw
rUDRQ3ISkIHGuRmHvvy3e+GgppAdKqFO92lFqsPUBQgxm4cnSZn6ZnKScayu9ArzHbP03C7GtfOA
A5kqHhiriQRgk6m3oF0uB7kGpM2Y/KlXXlt0WpvMNKs3y8/Ucwq8dJ+BsLfMqo/zxF19AFWsjbVH
na6/T244pCojMYVYSOW3sXFs9zN0gGW8dxy/Dte1VJjvTwUzOuNYNe9Mf5xGhjPMZBiNhEPrRTd4
O8BX5HIlRsIUFBLdH4ZlVQgy2HuMgqMT6pc3R0oK4asg1t12DFVMNcpBVr4thKILeFhEmjpZzAW/
Lz0EJeHLlEJKcd4fKQaTvZB1ACAGloqx0JaEAyO72+2HF/PYLE77q2frmToIMnf/srCVGvysVdMw
ROXmo1eKpuAKwHO+wsDctTf30+IqGg4pZFz/Q4HhHLY+uZNbxvYtL4WoQxO4u08cdzut8YwLgXK3
816CgluT6S8dkvHzL4ABObg3KXraRGWIIbXHJA8UDjShVdDF0sqM5kdzHWsj0rKvyAUDcgb7tvCV
S0gFCaLjxB2oHt62Azr8QevO1IFbG7e0fpOM/mxHzVdAq7G3eW29fJw05vvtxlGy+tEFyRb/ibZU
U11eYCT1FnagV7ANqFQpOuWe6sgx8a9Wp99r/h09Wjbu1tSLB6ltp+ahjruL6FDQ828zf8ftkQQb
JFh4DDasAaAahyQ659sX/BBweK7bOAUboKz4lQXQ5bQzJIMVZTNi9urw997evXdF3/q8BWDMP1kk
g9iXqXTvqIn6YfI6jcN84ZWZ/XFXgZ/SFWfHaaETufd0/1Bz4nmNo980JF3XEECzZh/7QYNZv5zu
K0bLyzGu9ZfyInSLuQeJrDTmBOhw/N24Z2QOmxNKzOReQxiByPdXx49aMkxZMkyQ/w1oy73z4S8v
yA8KeR6QqTTfueOLMp8ZLa6e6USUJxbkxJQI+3rCb+J18whRALX0vwut/tRJTsimEFnXYVTXB4aO
lduglvcOFOnQU5w04gQY7oYm2BfIx8e8cwKRQ3sDbfG1YUtU/L2GkWAIz0yWMmALoZZ8vccoeLyB
hGzfCq+lF8G0Qu1d55k1FyopTwNJNBpc+elxwc5lrZIbxL6UBlQ2Lm9PQZTtfCy6tW3+NheyJKTt
r9DF8B1lg72egxSrkicCs4IYVFAcXK4hRhLW6Vyt+TlrTh955QBlDWq2YMHzhTqDsXwdWx/k5S5N
0xvXzP3nrIIWwhAivFjk4p9P/dYyfaViz1tgyDC+CKOD+9qhdpxUEl4EwiUIDYy//OuMT+i5lRjG
D0OockCmbIT4I9nbWGCrF5SaTsE4LO9ZrGs6myD35TOrmSu4aynbDVjU0Zt55b++9RqX1jpWQYrV
gJgZTLvxJ+9ciABpVdkmLh56bUqkcVx5VHb+M0uSbN/n4dmPHPWZaB0S6jiO1n6kwHJnZ9R5QdlI
0gvUWEiMCxpAjtVIyps2M1kZxhmlPr2y88FImtg6EIaaEl4E+yvxPEoiyViskBQHmD8PmCkb5E90
8249ayBWuxOomz2SW+sb2uIWBqTP5t2iWeeUDrEu0AounA2M0ZykqjPTKEH4y+r6aflhj/XE2wqZ
LDfe8JeYnDMYXvr4XGXJ/zkYifIFWwupKY/fxqJW29e//fpHAnUs5Ve3x/+ceO5pBjDeZUeDyX84
GzjkQO3O5QXRKUffutOWPijl+snXPXc+JULe8sX4RiHH2qJshWHprJx7vJgcvwQ2s2LrtLz86hQZ
oJ5OfSl3EYol6+vVcNO+I4hUUf/BxjL3DFUr03w+2kmIw1v1ErInLmMM1ksgONsh1+ZvXs/oxQpV
JamEMgwzYcDQtWJqiz1A4wp2tWt57Xz6SiZM/yJO7rav3W+YQYeZBHZ3w1ZjeAnG8E1gnj9CbYY+
71j5qg3/6WGmMYmd/jmt9Yl93JBzRpOYidfgTaIietrf3SvKVmWa0Q2xSzWmvGohKTkHexnY+YgW
Pf1zkZmlTHciOrKtRnM9XsoGkPdDhF9PM2jDkYN9KKKvfK5nhiupqrtWinwqBqCw5mxpYGPx62Tw
NlJYkgfwmdFn/jKA2oLdL7sCjs4N3m6fQf5+EhW6o5ZhwG11qhAqD6APZkHYz2ptiS39sIlJNAYI
ApGL01Iog7b8CNdBoXPYhvIN1+qrhLr5uug+3+zHrnUv1xfsG+9tV4cmpGJQjSaLcjJa3azxu90D
0KchkQFPdrDPDeUe6UwzJbf75e/gxKamtRDNDkKoI9SPdY9/Xe5QK8HH5+Bbu5BWHhN9Tvn46ylM
GOVB7TI4U3Vc7bgQ4SGf8DrAIVF1TubjkydjvlmQQ8V1oyLScZt4uJrAF3MgwlE4qsi70ySH4Y9O
8kkP3DiNmhpqExtBsZ7ch1qyw9qIZsxyqJ7uYEUJBd4kr29JfuKNnP1PeOQuks9waPy9fsbGD/iQ
ZmAF982VwKIUmKc6G61qlq18Ctm3kTZyW+sUvIlt37qgYtbACkGUo/FJ+h14zkpY7DAiS7KMw7tv
iwfylXoIM8BX0xFCWDVJH3j+C0QXKyjxbM0eWGA1LNtEwQdI0+zJj0nkteWNfeGUhLuF2uZROWcZ
wPE7ssWutnbGknlF/guchxYYJI4X1HbFAOaOYKTF3hyI/lTfp3eZrd/GI9hKhkNgH/j+BigxuxhA
1zIUeEj87pELTU+VEiA0woPdxg7Ilo0bupyhGlPFa9AdT4JMbW+XJNh/v377iK7Ww/gHb6WL08/l
0iE9nqj6X6LE9EOXRLWHFwnUbx+hE56Js2mILn7xAAAuo5Rtd6FQgKtdvDQ/VKEO928NJUqMy1yO
aGt9m0raCUlfGiwkBLmfwE4LQ6ZmuhAVbcTMzH8InvB0IloA0ejfh1aLNQLdef3mYKDxo1llIuyk
0xGiwukxZ3Lm+Fg7LdeM75RukDkrTeYHLTd8980BiFrdY17jEO+mnTLG5to50zdiWlKbnLRAwtqm
PUQoh4CitE1mR1yCTHQ0bXS3FAvrPz1EZXh3KSMTV5iQqeGDVUan2HV+5buFVC7rpctTUDp6/DRe
BoPlcZcAUnDhcXtS1XbJoTtsyn6o55984YiSmE1vo1stpvVYD86GW8IZN2ceZXCzqocb9fny21ik
H4BqP388uehYewZ7Vip7g9GKoGIDDyd4uW2cDCufYWvRg4/TQOkv8xuPdS/NcpQtN/S58aKg/8+p
2mYIE1nqIB7f9AB/vL6A/u3kmvQ8iDPY0yOb/WXmEAjVSSF6SPDRf4ddwv4h6IvNkqVVf9i/rC0N
Qucum20W1o8XcTzt8BJE3megT4dRhSkSe+j/ZKdb3i+AUZgRvA7ZhjYOOhu5cBH9/JAFMuthLVEA
U9lc3/dVk2fSJd/KjYrOB6V6QPKyxcqyYHjzREe9FRkIsK+YPefz5FjAKi1u2acrek3yQ3WCs4aO
nSrTML+CFx91kIk/hyFpOu8+Z432PPlDrDGHJvbvh8vDv2FaX80jKbGweXho0IuCbkJ+wL3F+E2v
CAM9bS/x0aCXI5DrKIWbK7eopaPNkdTZQPkFjxKVTqn/ZO7x2o7Ged0QehHJ5Z/buwBeFoa69/+G
9hxKplAEDiLmmUKnPdq2eKw6bBIkZrjPKLmTtmwAJP3SR3EUNkFX02KD4qIIIgm4NX9dc5ZekU25
PM4MaoWfnHbAJIgQWjRiYxT67XWMnvdEKCRw21MryZ48TK8WwsmxyDBCC7ZqZegZhhTGXqxxE9h3
U1s4cRA+oRO5fnQhAAtTiNvm/1YtrlFqVHtoxW3teUZ3o3UymT6QODh7x3KNOXK7XvJg0LMcn+Yc
w+Yd9ByZefgtsyvVmaMxEQby6XgVPqVto44UXPvQwJtoEkcW/IU0U1ME+PgG137XuZXjorGvBSq2
QA1lidMg5s9VOmclv2kw2GVh5XEVLylKS6CK6bu56nn7cll7DYaTrxX16QSSZm4R8uhmaI1A83x+
sV4VLkgM3/30Iwn49WlepKQNTNpPcCumPUNBB+sH2P/IxUfnOVF1VLd221Pye/T9oO/vuE+pYYPF
pJ97IwPQ6UqwlOiE3Ib9wlnE+sXVfpejyDnAw0Ff9BmOlTU+z+4PW8URz+37J2mf1vYrmnTepSJZ
lacAwe5D+4H/wUoO0TqfVH5ZFC71yzrwDdbvPvE9hiKzxIg4uCgsXlx34hMo6rccXTWSpigDbF25
xUtpn9RyYT8jSIWToTP4zuGT2eRt6yrWXoXJ9iIeKBFNgy0Jo7fl3jK77nvg9H22ndVEQDiq37e5
Znj5JvIOqr42/UWdDFvYfysYFV6sNjmUg8fadd+i1LeuzkIL6e2zu04d/qfWYzNp5JADRkGy1xaJ
WXTXhpM9L7rz06DwvrfQ7Fh/habHp0IgF9hlykPwP0Exc9F5/xktMVRn+Cb1dobpxSReQV7bnir8
UZqfv9I6QGimc8GjxgUPLdy1/uzYu/uNqzjNAhIc2hsi3Ds9W8cqU8JF+dfL5/KnzFvEu4qGjE1a
wu8al3pa8YFEELI81vHxiafmGVZ/Koy4JGAjCF64y2ef7z4NCYWDOjsVLmQd70Zddz03P3ecZ66C
IJ+BG6WpQ0Ol6Uci5oAGieQGCLHbW9ygDDDXxthcwXmJjCD2A2+l268NR93eLz41tdMVpSS/SDWf
v2PxNM6VYh1E82bcy0F0Q3ytrxnCcmm7r9biNGHtgesYzGo1c6InshrAdboBW4FHAfsyc2x21wNU
2dARNlv99f0EXeS+Z1B0nnYti6q/WJ7XF4/3OwaCXvfCilMEgOyng91eKAiJxQ93H18O1XpTF61q
7gWHZ3DQgE39znxtNJOyG/onEfAP0GqQofHCeD8pIadKmPRtb7AMNO3jV4mbmvAiZv9r3+av321V
zR9nIsNh26Atucx0K9PLWMVSl9bGFKN80CmchfqszpXUt7xbfBvTNjNp8yI/4HvlVO/kVujrP+Ai
zhpwO9rvd4yneYkD7ySTMl33uHA06ln5m2lHBdQsfxFz6YPt91WyZtbppV9qMAm5K/cgZGCNJucf
weqS94LxeED7pftKUQloXxOs8FHYcCt9N1o9khujudgmUqOl166Sb1KR0dAxS8WNhEDzaIhgiNJq
LmP+kkEi521x/A/jYKrdK5CdUmIqGSKxsyMrwI3AM4F2apPA1vqr+93H4dO/N6GIpanVDG+egX9s
l3IOtkWWvmdgQPAZRO9KchPuEJz97SzFhzdGxlAcOecBAvgcFc58iw4+vxteE8Lp3MStbt+8GkM/
0NMJyrzbXc2xr1w3a3uHG9FZjnMyEpBKpXjQYHFZwSxLUhwklElxoQQDuxlxqZjk10G5N8C41kHL
qqMG8aac7uwT7F4XWrtgGnwznTfapf5fZZX+eM+A2Zz1gH9++957rR60SOHZn1xdYRZbH3L/KfSP
Zcgn1Y6GdByWXnpG7DCnSHy7OGIJRkgcXuKQxnXPR3x8CJs5AR4mreQQmS4kNSHkuhdlTQcrzhwg
Bb3RNczzSXbdLq8jdMTV2JdBa8h92J/WfTmdSSsW/VOqsI7I8tMs9TVm//+UgpPSX7A3w0NJKhgL
PjhKRD6TSlikGySa3FFRKa3WpvUXMWqlCmNtejEqbGjEWL3ckH31SR7BLufDavtqGvMXS7E1je9k
fATFOGOD2ptNKDHLDnoC9QjXLGXTdbLsxHFzKJsX1d3Uk7eOXEeqRZi20frM0ZPnFahDgjISGcIP
jIEFrEEe+LSjK9MxFfG2z7fUjq5kAL3McOXCy2j2FCX8ENefIQDeBmuTADkgfMNntvpwvxiqfmq8
xmVVrUrwc+90+SpW5/2Sxc4xH4nzrlLmQ3U1pecLJjtC9ctW/HIHMEAWJJoLBBMiETiVxmFV2oCT
0FovdV0AZKxIQogk2Yt3asXtxk/MFpZPfukgF8szCBgGjc7hY8hTLTBwHzuMAXS8nJ/A3PjrIedE
HfRP/ac1CPO0A6/JzsQETIaP+qWT6IuZfcUxN31/NiRZyOCe6/QcWQPIU0f326AwO4U+vTBu6+9m
7Cn5bsgA7w1MykyMjxdVWBUnCXOaN6NrKBYPO2rkLO9tCAsew3U7hwH3yJV1ZtwvEgO3PJ+5kTTq
QL638BYeVosbkXIl2QXUQqd1cKNoFh08+rpVkhlQ6ciJ8E6nlllvBlmGkreDBdCaMpKlQbWEclLB
PIwb+DwpqIwopklM2YuGl9c2lpbAAMlXvTWS4p6iOsEHJzbYcJ3ZkE4ZdUOl3a5jA/Lb5wuUqXlG
O7FXsi/ZWI2KDlguiBi2VOxYMhytp3vFquM1GkgzxWqzuUKidlhAvo9zfPfvw3o5c1C7cjb4Zi9W
3cd7WEeLTEI1Oaj9llyCPBshlnXKq/NM0b3NweYMga4qE66+oy274t3d/AY3ZPsaATFmJ3oB5M+y
5u0Gdkr/2ybVINwYQTVNwYcLZJ0Y3jX8bEHjw2cXY6qnB+0/jxYLYbZqn0zjT4t7WSfGEVMRDpAx
8IKjpzQhfT6uKkEzwQsMvjFMKcAVrSi2suMx7VBjm8oIekS9IJ/ZbqQ6lOoQeIcwGoQCezJaPptp
t97UmrrfR3h8jVinqtJJF7MeqWM+ZGWz5yGFUBgX8Tsjkffj7J3CpYOkD1yi3klZuhYmmTa01W4q
fBllAGKlVh4CBm7FLO6jrC8P1hi87mWVB2JS6/MgUoxDfFUydpUiCDX9NZc8AVZXj9+Zn6UKPjb3
5m1AxC4nxZvk3NGbTSiotHogPOCMiTfSQwnjsl0t0Puq5eGd1pTSN3j5Enhc4y5KnRgdAIQ0RhVg
CElMAuvjp3NHmcp6lZCkIcpUl44ftqcXj8xF3kSs6xXyXrKsT7NQggQ8MSxALiCG61mTkd6TNqDa
fBAEiJH9SBwLKR5WToUkiYggTMb5b15Y3flfvSmLSCp4xg0n1HukUceeMZDPCdkHdnDMe4aEBna2
5nGfM0Q+kPh2OfBmgABZn0h0hhxaYEBpP0Qjk4dwArtNir6aUHYPmbTtsizNVasYorDixdHnnGnI
KAUZtjLoL3KQxNAkE444GodtR93HfswG8ZNykl5mfdOa8THDaKTudjSBW09rHlSLfdDJybyrjSTR
0qTCN7sfGxM+zxZEmaSTWGY3pwI7zkQl6LrmK2PwjNyZAgldSA2m/FJpbs5raxhL6XpmtIGehvho
dii+tTFRPyv6OSNb6yyHxI6Udlv150fV6oRDBjzd/o4W9D/1ZQ2kS9Q5KDCTeAiELKdAsj+T/xGn
gmhani+Tb9BSbeT9Os0pdx1NNE8x3Z179oJJtb+svqr6zkqlsLYQshgEmJutB0oWR9uuC2Scjx7v
RcJ8ALg1YG6/GFZT32TKuPr6AMi3nsRzyZ7cDOyG+IKe/X4f172Nt43KaS54Pp+BAJvCuQJd4mGt
TrEOXUq/TEhr9aQzB2z5ddydU54Kn2xA3Gf6SeDECW+ods/UzdeXOPkNlgUfamsky8qMH0fVKN+F
H5Z2/rydq8vrZs7TfB9cFhvEyG/5SagRjpT0Cs1066II8Aqdyn7fJ4zScv6/FIuuVLM9d7gQOV+W
3rKC/t7pygvZ66bzPrcO8YfAqP+EHuM+Wo3I11GxV1sUfLHr57+NQvnUWWTiF6BZXPKWBB2cOKfu
CMDwK3YaPgPeaYnSAfK7ynPtgJV3wBFYISfI2Z/MaYBvxoGaaJziLBmLamsjXyH980MypyQNmK2W
eVp+NKw+ilaueQ50U8XBWyHKIY6S9N6rflhgIHmbaL4IpI52ogB85S+mVOD1PLEF88nscugGGpEh
zrcbZFxfHyGOqFqc5kltA61nyfpXZfCUHGaHR9khhKGFh//Xocofcdq9ZQfJeWqHuoc4Twytabz8
P2q27N4erLCVJyhVsO3lTkVbhrA8vHVq4IRlGgjEGVR/xwFxNtWfFwEPfuFGnJActoP76oadYznU
zWKio99RqIDc5ik9IYFQq4TtAfqgxIhKwiW3VarQMIbiTfP+6OKwhkfxrDuFVNv+nRJbGtXiZMxr
mhKqpJWC/VDHHE55pUSaF9NlW1PXW6m/ChgnDeclcxtlf3hs/RyLZ4JkhYfVDcmH+r4jGW1yC8aO
Pdimg5RKbBjYBiZgIx21SWiRO/T5WaOrLEd+TANcPZ341dRqg5BtN7XqZLSn9d1k5U5aiaEl6BJr
zhDMW+WdrGTSZtAfxNcdzywUPnr/Ae297Hxk3+bRp2nQXdDejMxg7Wy//JtSTbO3W3bkPZ0A4bcW
mR9LivbGTvB6YMU2R37x3nliU9u7vTQHLZXEB57ccPp7i5zrCa3AGA3zu70pC0hR+62AUht/vBZK
gtxzbM2NHfw0GIPIJviAv64iyGeOzVycRsX9d2HwHtnZJrq/OPYhdJvIa4qh8VxcHvHt5kqCSHVJ
V4//T8mEqWymegv6O4rtgWToJjSRhXqrOCODWF693ZEERA93tbpZTq1mJ/rKQnGJrOxrPruK3AGp
fMBIKTSxS98v88+/1/1YlDQ74On+f1bLyB9DqkXJqaMZpNuIDn8LFDocj3AavHRDUKAl5ZnDEW8j
s0McaZGUiAyIbK9Ocgg+IOgPMiVtdJeGBZmtD6/1c6AfpaIOs1YLLr2pzcIgbBMg6BMwdcuQ4PVe
1idOVI32HUbXPIcebBuPKv2emuo6kVtHdrzkaaU2xZTX9bammubIYEIdQEWzVC5Kx9qjPsTjOI+2
rQH1Lv3gsugB48wRFro9MHDIxDaxzHGeZkvYKKAPXyQxhuWHtGWuZ0yGzzB5NRfCxSP+b3pUksb/
avVMKhv1UiO9VHAy+MI53v+5yNS5W4bXHoX7m8wzCFnbBiO4qOqsFs2maNUy+vV9WrALAIRfu4F0
z9vYhcC670XFvhv79sNlLyGZS3wzeLgSZqWaE1C/HFPzglXl3oSDbwcjc4MLX08J18k3x+p6Qvvu
sHXsspQiMNOURf9rpC1q+O9+RtPT0b4Fv8wzpZUmeXU7zGn7CNqSU+91wyg4E73n88E9Q0q7Wt87
mu1eXlmvXVYfhiRwB6hyd8E1rC2mZsdLuoi/cm25JOxGcSnDmZWUwb6mg6C5TGdreoYEq06H23VE
mrK5Hg1pxL3GNIDOY729OPr5ipnENAMppiOl4DzPMBXSrLVtQ4ahxHfQ9H0ohFS1BoqJKLOSmEoP
JlBWajs5NteR7avnieh7THql2YuKV4Wuic78FEFHfdFGmZrjLIWPzBUKLkxX8VfFTMVvOIxD3c81
vDst9vwCM8vVAWxhIcmS67JTRWCL/ZIHkz6TaX8ajImmwrvE6TxukbMZ2oZ/xGi1KUFt3HjzVugs
szHICJBLpGTDP4rkO7NEVq582U5xLbIxfrYDQW+sYaIUEWv6/tbNXbHeTQGkTVY/jgsSz8JGcmhR
wypXZs+vXifkcPZnelBXaByBp5dJ8VKL7N1hnsN/ezFfvKwi3jgA4xXolurytBiVcM/9BRRwmeBy
noa9flkgn/jK3P60e4ki9tuug79rRaB907Mee2NZFQTxyfCILps1MBHg/dmDP8v9/C37JHCyjjj5
DjQnL+5H7s5ebL07Hyn7Mo3pKLGzD4jMrEciXnsgtYpL7jOFrzRvqW6rSg4OJ1f/DKIvS7O1YQhy
jhcKPHzgWzhzh5nfE1hirkeFlqkimZHkLHhJEbk2F16kAictd1rabElVVZedJqqC1BBBoqtGL/Ma
kmbcCM1c/nCKfag6WYhXzvLNqUVPL35XXp6cY/Cjm5jtz1UfxHDJSvtGsbEN1ia9HjD/DPEDfjXP
QAdX5wrZF+J7zWPXtbhX+DVof9hROPjuy/26vqhzhzpqzvfImy9f9CTfeu5+rGLqJV0K9XRvRQn+
lNMJk9Oy+BXEIz6/UuvL219+PkG22Wx/Z+IFSpsq4Vnk7jSm4Ltb771VCVLlGxVCKJqV14tn+e1a
xF3GM0q07xE4my2LwbMIVmQwxYlHnlW5oCMy8yH/3WQ1gj0Zm5PN5vCyZDrNLeViTyv1r5jFWHkg
lGr3Z4cChSby6S/vpt8k1na+dbg6vQKrEpuP1JKugonI6OEVbzaIIcZM+8PSN5uS7ZlQ3luEJdGu
+D0YDuFkJI/sGwvKPZrYXOGHSGwrrMdtcgwKAEYyHAG4UdktfiIbAH+2NYTfn4E0KTYBTQOUcHFu
XVcNCxYDOU7miVICbqQNODP6CAHuQX7FFTpiRVJQXSZBPXGQ8YUXsEkVS9kOUhzh0JUF7Juwd4z1
9BFtN6mZxK6KJKUXeP7J7fPmZNpfsgQJkjhTI/LSWP5SCQds9qKQzSGjH0NFl/I8R4CO2PJNpi6G
8CIWs+Snuz0HZL8y7cWsURmTFF0lBTKVNj9rIKzX0eFUkDWIlGHBjTa0Oi+IHoGaxgShCNfipYRe
qEwZ2rfAYUbreNM789+k+y5K06eNH+P8eBzCxw3gbnU5E6Evs93x0iheHxcqqk3gkU7JBC+jrjXp
AujgIXqAXWutu5ZCcMP0cdJAv5Iq9LFGbbHSnMyTndXnRTbDeqpqvBg4QUK3amrupTYg7n49Cl8V
cux2K0kMAw1Y5BBot3lgRLcXQKy5nasDsoCskmCW7E+Y4i9UOSyfO/eefNlIb38QiXAITMbVcNjQ
3KkYLFe0L5Wdc6RMlCJ8Q4Wb19KgVgXWza/7c8xq3tLWJPbpPV6dXF+wVnULt5ufct/h3nb4ih7f
aOOF4ebHUw+EEkY0/llGVH6OzLoZcniImnPPFNoTOPoP8+6+jfVHqtZsnbea6LOHLr2hZ3hRk9J7
41CqyKA1dU+109PQLhAnQUgLzR/IIMhUlGB9rBKwCtjJ0R7nd9fZKHb62CXbQQGxfs+ztCrMsoZj
geGHqJCb4hYwTct3IufmTRpPuzTgY4kLjQq13RIA5fmX9Sic4CDl+gcEVl+vHSTxMgYxgEtx65LG
D1hecBp7v7Q++KFSucjdjFyXrvXHz3cgh6iEKC1TnjSlQVeG0nhxL9xU/zvLdMfTnqGt/dVcEL/4
CZL0uGjSiea946Cd4VYzDhowYb63PRcAQf5aS48vTS6s7OhozwKZD7qfoRjTAhlq+a04tKgDRj/W
YqnQ6ZAzdOGKj4MygkQvstUJ2WGUmwLwzadrSjPCqPuSC42ITvtDfOrv30UC4PsUPAwpP4JlAM85
Saw3EjayyYFLqVYqM6Xg2j8lzWeTueInSKCznRWyfwvTdkdDP79Ke20jwgexJ23fFW9zb5skg4h3
lIO4QrxJanzSdXARRGX5slRv3M6fmUFW1+ttt/2FN7rj1LU/w8cabFiF3WI5YIng4ffnFlXYieQe
PRNUN6fhY3TXoO0DXGBqT/9COriDKlZe4t1CBAxicWJ0jCQPTYQIWUU0zyoN/3IZGeE/OEqVmxlA
CVxadxTazS33Om+1GSdHI1gSMlDYyf0LAJCpbxmms3tK/uHZLwYHfRvfGtDZ/OnwZT3VzffB1jR0
JWdJ8pgHK81VX+EO94HSaSLy1cnq201SZPkB1vhdWge3peZ/7ay5DeQXzRipVaq3j0rmbTzl+CVm
FjRegOiIqIgF0jpJXvGDy9Oc+dbtq47KBCy1A0TYzU8MGcOwugVcA/h9vK9fkahM447MFV1Xobev
FN+LT/2E4aSPfkHqpQ/vCHNPeLMCLheXZhmX49Zr+B8+vutQiofGvIB13KQog405i7Aqa6ac1ET3
WrzzJeHnZJj8ycZ7HusGR8qtPfiT7HcEqkl7B5llvkxw/O/AwR/NI/QDZR+6kLBiINZIic5817/P
+N8iqb+Dr1XNVsUS/Vjjq1vetMDLwEAiXX8ByQYHMFT5PkTEY3fY63iU3JZ7cu5dmVcwXTUIkUQF
qfa6dYgdwhwJsNRjDgRo+G0chPY15OCk3uvUN6CYDHEvspAxg+esclSdxqItugRuORgso+1w/nKv
1m/lcf4+R1lxisysmAdRMs7jPwjASa6+DS4NXf3JcTasC2paK4SZby+39U0ke9I7+8jFDchXt2qb
YuR/bMQQQmwfpFq8lB4YzEW7SQsa8txJ4Um8t7B/6F1eBh0AT3GwTSRk+sZF4gYfzNvCn3jFbj/c
18qQzgaWZgReRyRKifoApUwKLpfnfcaajNqteLVpW4p1ks12wskHnIRUGX4ygOPiLOejUwJVTldx
S74Ni2cLLWc0IS7kNp6H80wvpBC8Da4FhWTNXFsVVQRQrPjL7re6hPmiyXEp+WXv/XBxJvDo83BT
dcaT+Aym8RqhYv293L/J7fxO5MdHEUs8SMefdScbV8a1Hxl3pp6EZx0teoqy+wfN0Lef15VG9ZBh
Z8AOqLborvzwsHkhei3KieSYjUtpbXbw2tMjrnNg5jRfGzCyHLGVFHf6ktzjbSBXNOWsIARNHCSc
d5rss9pR7B1R6gQPy5NRMHwiIbUW/Iza9fLmsG2Q42MrUHhE5qlSoDv3MH2Rw5AozlASfTNODkmZ
7zSpqEO5cczlWFiMy43NhefjeuqcHPK2ixprkf0QAfUc+z+xz0K/eJwm6ZNg868/zqyM52nAL8hm
vhdohxfBoIo+f+SD4SGGWM5LJKGL5DzfiRNSmjfj3JugDMsiTx9uSMzBHWUjLtYRg3raRAcTJGwK
ldNfPbaxpz5m2vztQlKv1aDArhAvgBCcLvp8/q0cwIdNzuevWVh8mPMn7zovwEGu2wuJWWAt8IEl
KCHlSxqdqwhFHQDS6EIsakthD2QEvExqovnLZqpK522VKfbxlquRElBhi64ascWHIcTQDH06o/6j
rlOhJBDKuTwWGY+IgM0MQqd/0OdvDNklfo/GStT5f8EfiV8fuU8ql2CgvTEFBN8wp1BK5cQKxOHR
6DSMKOlgBe6ZdkyiyVhqtrLTzkze1t09VnpnGwUyUlUvWpoYjkHsouWLWBS/LIUHoQ/aNT4DiEL8
JjcQ9RGWOD+Lq1ConFWzEwH4ViK/7fQ9VvY12kchrDa+IqbcSeGpM5IF1z+oUBCtiItKoE8X8YX5
NiKbM2dGx7f6GTqto579D7DjHSnenGmwRt5izrsWSbBmYxbHHedG9TCGFjPJPz0qF+nPF3AMcJac
IB1xFkVNL1o3rnlvR/hKGssMw18p1sVFmJs5QNfOlviPUDylRkyDu6558LGMjgNgCc2Fyu2s6tH0
zwmjFGbyDyRlufommSHLy4WAwwNaH7V8MLQBi9Wzepq1807lLFhb9PPuy1edBcn8/98XykXD38eT
V+z88mGTFjiTAC/h7qjVw3jUsenpgl3xKHeR2XxIs2pfHHyrvrcR9ThYCj166Pe50TrEHheIavIL
/pivkfYpfbhL+VhAHG8z7ltdzS59H8bEy8oJ7OVxYvzJzW0+di7Xy9ogj0M+C0cxnNEqGh9me32F
AhKg4+1s71bqhVBgZK0EVW+v1C9UhgRjozPFugnG481KVbxsvBzToRLvjuSg+27DE1pvaKK6nEdW
Vv8LsiH9mP5ZMaJWzMLjvU6xQ4AMLH3QA34toX8s7bQd/p3Y5GJ1h5Ln2O/bgOJiFvKW8npmdLjB
/Vb3wGe0lqFkbMUcGODWpR3hX494nO6KH8LsCZhbCOuZNtrPfbQuUL4rVUsjJdG2zR8V9XxYj1/A
KPV7mS9qBnCgRQUyPrD8/OWqWl7pqGj3chAI4dVJ3ICPWuEELCrjowBeKy2GsjOSnea9e6NlGOJV
zUtzjQr0TTXjOQWKqw12lOp9Jhj4RRw+SsoV5PpCfXQ56jrnoTKjegOmo4GaXlFWLzBA8CAMXnNL
i2PKwGBVsUxmrRDIMIpBEeH26VUMIwY+oLWBlQaQ0yJtXGRomAm8mlor5vevizJmuRNB6AR0h+Bq
07bDoPd4rQ5QrcdW//6UXSnOthhm+h99t/c9N6lZ5pP0eUqEFN9M/rO1ybCUVhhb11dbToJg0g3Z
OxrgNL/p4dZksFRGVJi6E8V9d9j6A4FnfU+HkiTfmcVO4Xw0HOt+xE/KMkWA3H62/I1ijMZpR+aj
QoE4DAPn6Vn7D/5UhAK1Piub0WKoREqgAlyrjRuH/91pzcqdMWcdmgIg0bOZTgHJ4iC9yatktqHK
xqHaQy7eGUdLbsvS0HFP3H/ZeDGWHc5XcteCJHbjenizyb1Mfhb44BdXlxBWEfLGWx4b0/0PrSrc
t2Q+lvEV3QKAua0AY2wkBmsOMpWEkN0VesDq9tUMgkwQKPvgYJQB8AZ6x/RXu9E/31X3jP/S5wfw
I63DAJB9bYugHYfU2i4JtOdOwVMLzV4e/Pexu+YSxZkP5CE1pOsQAD467R+lqdLMjjfbXrJV2re3
2U1FLr6yFeOtspVzN+P3UM4dkYeLUBGRMEhE4uFAHwzn9SblYK06IloyZCA7KGyLCca1yRPDaE/s
/DaKOEw8z+KrDefRQhgVZBvEWs2/DA9hVujLUsRaYJrwwX3vmaMBdfWHkpsf1ibjSjAVeNFmJJeC
78+Uzku3VhFxFJ5LR2QAQTJxQbDRhkc1soP0t3Aa0Ngs1hvoZGiV9yPAZHuoptfq4dzzDVcAsQXS
SDG2qgV9tG4FtbLEYaDOyxTfyW7Y0Lv4/cjpYhC9o3k1Un064fcjagfp8xJs/8R/9j9cr/GNUzxM
+XLVIHfqcZo+WJXaNRKWsS2cjWK2lCE4dHHaDB7vG0SCK5zyBgShM+aPKK73yzNSRSdkccDBpYeC
g2f2zF/K6Uul4v2y1hVp3RvyXrb0WJVMXpJ8segtvf78LwQ+d56u6gJICaa+G1nhFnkjM5+CdSUh
q8C1dpRt2nnfCFkbhl8SEbDL1wccKMkjMQZ7aL3hrKUgAMq1Wn9B8C0U0KkIwqRvRYuG2bDhF4YO
PWBhVeV2gvgRsNW8ZQS3A5tYlr9puI4AVjlQTd1c8drjK1TxDXJZ8jUsn1pgQXcx/nOIvsGKoMC7
iYxtrTtRZ9SXx/t3mDlD5unFcHWwfAyLTwztru54Ng4pjQvqIDvWzz+BnnfIMsywlFOErL/ISFwx
UPWC5Q5MtwDytsRa5iQIRroMyU8X/8zQEgcFLvtkat8hcEUhM/DRNoS3UUS72MYS5tqfGvY0aL06
esnQealoLpB3FgXG1nT+4ET0Z79wd0Jj8daoWdRuplgMNT2CUGPf0KrD8PosQ5Dx7Ebv58FBu6GQ
TFb2SVC93q4T1xhwVjgIojAXaviT9na8yVjHfS5+IK7t9XNtnObJdwOJ9Utzzo6oyVjwb6li00Ad
iTm9+QKUirtp2Xqfn5eAEh5Wt1gJpBOh3hqbdw95a7JGXo8U16Z5+yjktH1gZLAcWfiO23X++P1d
gpkaCYP55qA4X7WX4IfMgIhvpF0Fglk4Tn97c3oNuRJ+opdNDaXb7kZRcUVOUfM8ZHQvBwOcquLT
NGDtoHIN3olu5dskHQSvfF+nKhYPLUt+Mi4MdD6BAf5VNQ722K+2AU46U1on/JdAgYQ6chR2HlvN
pHBfElwyX18C4DQEnX0cTeWhSoasW6LTJndfc0x7ZyzqAUAB7fGRj9M/t35z0t4OI4KuVJDjmtYv
nvc+gPLemuxSD1G4A7IekJOJ2RqqJQQhbqugH1MCrs3xjX0Uzu4MBD3osf9iXyOmLsg+tantQBP1
TsMH9NAcxXWyDj55Si+32z8/iDDyyjdw9yWjhHwWAAez/FRpH47NQkdO2R/MUF+1dM/KzuYgeoL+
aHqapIX/DLhPIUqvMvz5ZXmESkhoBnLTJ9WKGJA0hXj8ah37X5tUXxXv/2pVFE0K+ZS3Z1lQS5uR
THhid0qDlffF6bIodkJVcAbohf+tRXgs819kWbm+93h/xlvZ/yhCf6e3RDei1kz9TLr29yjapHCS
78HfybSEPCLNfCeNdI8pEUZZRm2Y8G3yag48WKP+ACrZBIgJenZySrhY5uNSdEE0bui7Qw16VyAR
0F3uSj5rUUIx/j9wiKQ1gNnv0SYeaJkHr69+8Pljh2ijTt1uLvmGKb2sJLf5R/GHxDDklUEoUYO5
HdOjmm3zIbRYAWqUG7bSIKOrRrTBTuTtVCo1SF2E9PSJTDa+xlpZdU9QD0HcBWTyNiWHHXDkGtCW
iuHgpQzV8JIDJc9aZ5Cjl0j2oxKEvGsIAYx/HVY8jOTE38jZS813xrAQCJpGfXUsa6FhBwYldl+g
AvvQIaD0d5xM9dfiLNItU0CzRUDPUKP+reZ4uAnH7em5C4SH0cWzNF44OBgzml4sRNw/DC2YFgUr
mfG3M7Fdv8tnA6NLX6K4J31Kckq9E7QY58YQhW0L/PdhhNxIpG36cwq+UTySqhqEFTKD66l7KHIs
qKfBBpd+LOOGpGNiwxNyuOQ79IJd1U5Hn9HmT2yauqJsGDTpfjSPb1R0BavrNKB87d31IpCfzf0g
6PKjZNWmaRmwmV61FvSEVKlGXrIMU8yt3lnc89lvfBbYW5QP4K4vJx3RDRO4eMKAR7vTCef2ywO1
cS0/NenYkpDV7JuuUi+DSWn/AmeFR8mmVJ8kUMaYYtOM9AAS2kouJAXNr/S0tEGYfovx5GwqcB6S
KbCy+JHGzmk2fwoELvt/MDHtcFLk4lewQ1u1ZUd9gSd3ghcFQFkDjuLx9wbxqdKyyeBvSGdhVjAe
qbzP7kE0/ib3C8kLCTJMLvq3FJuYPc/jzHHt/kQRXoY3bjOuR3E5L0ZjV+fw66uMjnvSYm2TtEkF
QjJROJHSbLj7GkaLKUSK+TPTJaaVW54RWaUZNomHnepQnQxrDfSJzBndhvC8MZuQ5gbYVmR418RZ
iRrvJX7GbuDW0bUjtoqHYPVpycfxehQV7KhVV6klaUHr+3hEafKizGa+KWihtntYMuqzJ8q7uVGW
qKsmSWmMGhR8aSf51gO6G+UDUfJAdLOaXScFfx2dpvO2ExKE2rYt5ceF8JH7xqr9YdgIfJXeueWU
UswdpPsSPEv4NsMie+uxfJ1OqeZGUT5ky51wC7ZzJnsmeC90ulix6ZCn3N1ezg4oNDAw15VmdsZ3
XoNqkMKuH81q6OtI3tAmRKPmUh4LsuEsVJCff8oHnhSaT+gmZBtGOSMJrmNj764yNSOcgwgu4+ei
BOMqPDhv/B8OITLv4xd7dh6s5l6cGc8/kRJM9L717N2cAd/6HoKX1IVQeBLaiBTVN8qWh+1Jlfdo
Zi63SB5QJaNnQzehxwUxsfK1hDv2tyYjbi6+VLIWMQ52VJ9O2UC2moKM16NR5VqKD6eKsKSuUguv
BClLY25C6ZVx8nXdraaCIgFOcfUaXtaq1NmXirUW6AYrHteE6s3cm6PqulxOB41IkyEYHU/QO+rt
BT/Q5ZgrdUJqufhgiD/QFC/2s9XYzYXdFhrLhLEKNx8s47HzLehnqxp+ksLTgsGfmUM5jPhqDMJm
duR55/Nogoz0E3IppWqTnkrwyndiHQifsgeS1RyIqB+BSqGrKYQdgJKNNH8fMtsMYNKDqjVJ757P
xzimj5n71oHqqeQb6XQj71IoKnVTliabF0utmKbZ3hnW4ZyND/Hd0w5a2HiD+67SI03H2bDA49vq
xupzGi2OhJrRF5U9mRm9t8tmXMMWYcXPiGLQ2URx4r2LAL6j/QZNgSp/NEhf2Hk5u0/pjkm7npzC
3AU9NNImPhwHPcBq+Wz+9aNRgi+Kwwia9FDWiAA9Qe5fxGyXcb/Ln8rpRUUOhinz3eM8gSx1MmVz
7WnfFSeCtTedHVP7K6YdLw6oN6XdTu48aaCV3/mJHV7Qewe1qDmdN3FoQJDEyfZO58ZB6wrSx2Z0
rVtn7ljwoVIwFxsJslg34vSoa5QMqbS9N5x6xXxzDZqaY5cg+OOJldqz/vb+xZcRdrlS5KHQ1u79
PMrJfk9LArxRHxnGI6FYzMjgN1/k75AzhNbRcbdDLYjb/EGVtsEfWAUmyQjata0/GHLpH1lm7H7X
4WJGHSaOcrV+zyRa6aLJkavM0KNvJMY33zDvVxaKjVAAlGogBR9ehTYFag689ajvExCbjW0wScAf
W9JO+0B7UYiO0/5V82ML41o1gm9fab/P20t85YPca/0EA/0GsH1kDUxs8SV/NOKikewkOEBBr7lt
BHUiw6wUtqTStOte7191PYMfN2XTiFCKrR3zErDSjXjiQXfXyrWaewBl24giIQawOQs7NQxa8Huh
N8Agf61BxuYiOMay2Nqcg6MLacyGTrkn6KvWzp6hlxAb1hkhN5rd9ZcZOziJ/vS/SE7XdpiuyXsD
tWl9GaRxA43sYgeSOOdwE8W2UYcDunFPJiTcLr9JkoP7OpNeYbzMARR3ZP1nLZ43OQrZX2tekVS3
CszYaKfTMK5+8OUgogiHHfg2nGhbQwUprEKNGQR2myHy7t5SCIN57RGwoJyvKs6TM/uRMGa1JI8x
3ZES1zqqwATTjcyFV78zo8G3OPM6MPszjuGBDSllkesN1Bk0wcXGdfeNZuPjK0OknYU95HA0rf5P
X0jKjkmlkCKMubE8CFM5RbWeBFC37zoKlcoilW51X5D6YsX+o4+2FAVYtDdrSbifjm7DOqzLIBf2
Dz3M3FXzBnT7vFb4+U3QcQPiFU8v2Km3QFO+87IzWrJOeuin9GcQ0fpnFuA6ldk9dUFrkeyZCdG6
aP29NKnFAFliNmWxJCG+ESqLxrCsphOPU/DRpKeReEqxoLwefC9RDbYgQT2TR0Nu4iO2nYrWYvRN
3d3WFNnB58Zvu3YUVozuXzFbCnfOlT+F6s9jBzhBmZ+NwLqnD9X1yb2IoYNlbSH1c1yCGc5OvJGw
9LMixOJhYoWdLWQhx/7IgeJUEAChyIXDtt1tO2y5ME0muwb0R3pZEjuhi8reMVs3hUUriozCOehv
RupiShkDTt8QhtqlX+MNd170P/ESKoshuCjLKOibUWw1XoO7pI54awJ0QimIT68qmdIqBt8Xpj87
OeSQLqnh9NVK5o2oIb52cg+ETCxXXePWMZfb6GB5ALTUkLxFExcNvzzIIpgTaE0+NBaL/zycK26D
pcOLox6BDbttDhYWKk/+yvJgB0O3RHXc9ytmHeNvcKlGz4ZVJy3IoTqJ33By3WNzgWqIy7Kw57Kr
5r6YNUqQLocDXSlhbXNljMOI0Wu/yjbMBMopxPLHObLWe9Ui0qAz/Pp87d8ij7aNI34Dbx9sQGIj
aJksxgZrnhL4JMy3R3uSofNt8clCDSuTRziHFVOxffck4CgZ1mUKFwx8Ic1ANeotweyU+fpDVx+S
m3E1m4Jtmh0TSIi65TLMeuPpU7rCrBThXF/OjOoLZnIilIut9frj1Yz/nAX3mt/8DqZTdzoMQ4qp
2w/Q+B6Qv8cDbV4qD1zObnTfvLnayqyBTQ3n4RU4bW6+EA0hXVFRTyA1O+BThdNUHo+zZVhYvZ7j
aDcNDDYEB5mf/lVGUdjLyZhwSv8vlP/sjoX1sitDiZGxZLp/zuLZqZKY/tVuOd4sCD1cVXjNgKIu
L7m84Clktro0u3blKu7ZWeMVab4Le3ZzNawkb3CJvFQsTAlyv8FHsu9Qn1CFoc7Ua3H1dzeqqp1Y
0UCI9Ah1M7d+u5bTnYGG51VzBPTIBau5Rv9X6JmNxB0FUc1WKPkkQP9hELVDXPPrUuAwhAlbY9uO
8xA0QA6lYM41PZFFXY6CIuR05+QU1URKKRdvUy6L8kO6fG3Qm/DT4QgkzNkTE4X7NpY73vOvvnEF
zOhhEAIkfCqGMdnDSO/rc7VMizVOXMZWoAgyrqTdarxWguHZspdwi6B1JYVUUyIW2rONJRSAdSaj
ezAXi0AUNuSWxgFD/DiKlxhBuzA5eShQL0xj75IVks82x9MIZKf9v9wxt/77D6vdrMyrD2PYVPKV
5gBYUJx3pDDlfTaxge8I/HqTQYIo47DT0j0SilGtzz7t6ZNSvHeZRfM6PZ2xhgApfCtAUcPk56uc
HrLWk9iE2VCnf0Wa3n75wh0VoB6HcdjoV76mLh+qJGxn7l93iFefPtUVIBuxY5KjzmVYEJvLL8dD
0hX8h0V61M8YdnX/LVlxdwaZ4dD6yGrzobgPCACEcTQcjPTh7o0wNTYBNlwX7Xx5937M2oFU3cr3
kdLgiIbEzwuv2RWEi2FWIydaSqUMNZzXTSbqnO3cTuT1u7TCph4ZY6CVGQlFmB1EwEI3aw9LdJIb
7JGTuQn6tI3YNEsRjHiY9Q3DnwN7q0BKe9qXqfAE39svQFSWQMKMx8QEMuEsrqx9jP2d/iIHgR7e
qOFaE+IR7ygBu1wffH9wVR7z2iJUXoatGl9t8iZ2hSN/4nYI69+dyhWVEvIT+BwWZRNC1GDxcp8Q
tdxV8naf/lFRSaFtdHg2eqXkBD3W/vG5FoJ2B9XbuVehUqzGd00xvJPd4LxXwgnrITOQe2Npqprj
guRUGeYroBHpRt1a4i8JciUPBvIi8t0/hcakgwmU8PCaHwLbphMTpPUctCqLW6+j4/eTo5Fy29Na
Y5YjSLdyWr+aMyNRBxKXC97ckkjo+uCLCkan+45HMekne9J+Cw0yTzwedZW++4W8JOG5KByPichb
RcZ7TMR0Q7dI/HDwaX9WNyWEEvi7ilaJboa4VfwlYxhRMMAXPDOzBSkzHVKPoa9eITp5MhxAp1Fd
qW1OswPw0IYTo5MqxoNjO89p3Ks3qj4zyf9Y1Npr+bhJagIxlSpdrRgm91E5xKDMuaLTcJ4vycEA
YYNCNUXtL6rj9Fc/Le0yEvWtzCyMToPUoBYvVzYxA0krUfL5eRfRxm+By2IEvOA/5X3cs/0+hszN
iqk7pazd/ngROUhvQqq0yd2YZLSYphgeseZSWyd+uRTEaDS0wp2z3tPFIWH0zl85AsqFZhcIvCim
JTsy54RvA7lQW3b6cEuTtG58zvn0dOWCtVN9f6Kq1T2hYJ3YqukpGtb+da74xiHbQfUKnNXGQwIu
wL8QB0gB6CEuMnkz5DKbyibbRBJ6Uew7Mr7v34xl4AFTZTYIVeCwLbDOwwCCjCpDYcBOEZ+ZROsy
E3ZD/JUf8Qf+jWFRrngIotom//nbx+qldKUhSpW5S6fRMWiPXAMJpFywVxLqlJEx2ktymJJS/qP6
KTX1lSkZv9kM5ct2oibeFefvmRMUj2oBWt3HPl9HnTkVlSczUmnuS5+YxbebCaOT/d5/nVTKDRdw
soDZchvHB0g9WPXIXxLtL0MMbAHdMPUKoMx8DzEW4duqq4OLauJdfoRTfB/dk2rehiRpHHOJIg3L
5InEHfYlUVdusJ6vpsP0I9d4JTfSJITNq20bS8UJ/0bzeYpvZP7yBHyltcSFONIMvypr51/k6l5C
rGJUKnKeLe1RRBUYRwr+ZRh2UGzCJVbcFcb4Bfqh1ce30rgmBAzG9HonDc2NSiw2MrWdUuUuLeDW
P2WshVSbcdVBPz5CHtZCT0g12n/7nwVtigfd0J6imBvNKBagDH6ikGVm84KEE5ClQqPgl2RaHTdL
Kchccgl/Y4a7RgjXyMxx9kzywGsTvBkW/1qsbPdMBYH5bqsG61s5K9/zVuQm1AaOfNRAVRoqA80w
sJh6PnkAIoq5ECNZmFbwgK7X7pHamVRpCrvMoInXBlsaAKPVtZINzELsfOYbvHl1Q8MKGAFXTClh
mlmAmgzTO11l2reLjRath/TUWKJaBkCZ67xejdXBanLWkZMhYhvYUGfZ/YMxtPqZSYITNl0Qr949
CQJBSL0iHSSeNV5/Xhm012Z7qzyTBhB4zBdHGOGuiZV3aAWgXeqlRTDHnPiYV2VVFitFTSJleNVE
5j4s/krM9cKn4FaVx/drOo45m8SLtPiY7o2UN74nQd84E/sJ3LAtsDeyyU+l7GW97BIHdLFE6OXn
XKBfsJxhrJUsZrtDF/ZHKloRphBrS+afER1xgX5yu/tVPeU5DLb6v5BY2jWk14bPoviHhHcsz/Qr
7XiqixFeygDVNIN1fZCx6r7VRTzl6gfRBypnPY1T/8GTJyhdZ8zdWnjGrMrDs4D3pCE5m4ECiNQe
Kdvjhv4dqBq5avDMSsJw64i6vkuUk+GyccGZkmhSbnc9uECqrFB7kG3W/SgQ0cHuPGC3v8sFbhP2
AcFaaJYCEUyyN4VhAZJtuQ8UZg9lSsH8pvfn0PpQBebAQdghsUY+9ho9STj0qDdd7dUCJdABUiQK
E1ahoFsCkGTyD/DEg226cll3mINYNnY9l8Ock/aS3uYTadtgK5wCNYosdjE2yKBC5HuSaTamGapE
TJv0Oerg5CYy34jnXI02lGF7X/S/z23IP9M8dLCQs+rnGkgUs7RC4aLZSpJsPtz+3gt31wGBBVV/
1RCG24B8oLii2E0tZi4GlgSp6NwOK/ibrC8WELkE9WwUrUZkSQb+m3WourpS6IgLSy2yHmtD+S6/
FyaqWOfkqf/7ToPp61PfKbAsCIV2DFhGcFEH/fjWVeZVk1J4EUgpr/YxvyE5ooy2f4tkIBNVkoI6
sn3V/Ho9JV6qwosjQk9JzZ46XYRTrYlGUZH0mq/Zl+Ja88dM364vcuvAOgYzAjnjNWciREan4zmh
Pq6hknuZwJW4YtBGGl3jPFoIwjlfKZDxmJBHtifXwumt24EqwtNh+9LdZpBhDGUu4e1E3sxON3ei
aPEFVDij6okSElVhNO6rS+A7Z9WTeTX61IcqODRkAGfGT+/Uc9y1ViyRIL4ZeFMZR3iLe/uz3moW
AUAsZ8pg0A1c3XiGzgvGN37JdatvcdSBCLuFaJRMNBeTfUV1cyR1kzWAfgFMN/Puc5CSLOwMTGcY
ttEUnjWM2MbXjdk26sheyEqPuw6/dKTtukj9+zFJv9oXnyN8rmEGJ/hS7Kh9Axv+wbsrd6X6ay0I
kEN7gdAAi+3xczMizasdIkR4QgHwYR0ZYPylegPnKmjp67vQ0hxmQfB9VdfL/6epsBo7DZj+N2NX
LdcWoiRDojyWgSLKrCLLK+vYlOSzm6i4/Jg9P31/t+GOzJVsdCJZVsX0lHChAeA1AOkOG9F8H4Ze
vxjbUlXuDVofIFnQ2Ap0HvC6Z0Z1hzS2q8UsfIOg0o7mwqWNNtX2ZR3QMly6xW5ZFVeaBarJhwYW
rKURpC70XGFFN2ttLzXe7t8W05JpimwQb+3wjWjbF67f+n43Nwl6Cf/HD8TDO0BME38YWHdMsshy
Fh+SUPLAFA5mUEzarRsMxX/HhtgJC/ZaFZL39xZsYVTg7teTpTUDnvEdSGNgX09SUWi9SMKwoKQL
eg5fg4jCs4H+t5AbNQHhpOitAvFcmaqNDfUejHr42yVEbzj7GDQAqonQeczGQyh1Pcy5dRuLF/sO
WcVyl4Q0qtxWMQ7zxtD1f2CLd8Cvf9vqaHMHo07PyAN5nx00mIhbbmLLey9qJjyHxI1x5h/bcMs8
NDiDEhmDz7vSoSf7dWaeIQWKYSVlESZijyKnFhbIlgLBHzvyoRlsbA1lToX/QoFkr5ihSTJyjkSE
o/I44MxRLvoaCIW9sy8Bgdq+gEmzvHP/c0ZJt7I9Guv8piU6nh0GK8nR1fjyMPPXbv2R/lPl8Ghz
MLpUliDnmQN3j2Y63zypu+Sc0o8eGaEwuEupVL5LzfTyE6g7bDv8if1CpiGhNVTcisfS4mJW0WoX
Cpn58K1ERFI2Q8Kr1uBHQpvGOlrpAstc7INPeZhiE+d6vS/Jq5Ra6fa1t2OU/aZChp5IURE3gYQb
9duRM78C8RrhI0y4gzN/YvnpDHL+PHFzhT/9/raFfhnrmu7iN3RFQPqEOu21UVrUvXd4+x2l/JYw
go1IvCHyECW5vLhohj+9+/3pFz/T2Bwyf4V8zZARe2+8EH+J00D9DbyJxxislaih5mxl+x1BxEQV
ngnvxdOUt8wwIukC4IFpR/WvdRRIPRDGZM6XLNO0WCY9YkoEk0mqa0pFM4Dd1ojkhkb0T1y95puC
Z9+m9nldv/C1TKED8LlyZrV1b3L7YodPXJQP8xbvq6OXHus3mX48E5tPzHzUUKwoZTaz1+XZyzcq
HKenvL4Kwf4XlO0kS3YeuW7YQWy0CWGFFXyjLnxXOKMf295uJsQpPSus+2yqGOirn5vHYP7li0CY
wQcSsMutvwdzyAG6SxkYxGF2L6QHaILXBlDG7sHntfavY5WE4aDLKzfSpub6zRM0iCSGP3McugMs
IwfhtTWbm3sZKYq1uE79ja8c6+tlCvilGLr7f/Gquk/trBMw96wU0TnCPtykWDC99tjA/ddRtsQh
dH25HF9sXGObPi2AaJAPfNLGumwfY2g/zzaHmq4df0SVICXjC/h0C9C4/mA8BDONDJNEhbqVa8x7
WAFhToM6YUg4gLosLD0a8MSTq4E6AKnfM+VCe3Zne2YhLCd7vusZ8NwrZhw+30L6W4z87eBWrZB6
XQGQeqJ++sx9cCF1AFhDl1R9JiD0XlX4SzsGS7bsvDFffaR9giKY1rC9Q4hjF89LRZesofWH2WWf
KVxk8YZUXUB7+DSdr49kh5smdkaRgz7lOFAwQGFbBqHyU3NLSNLp58D9354jMm1fiwAfD0VkSNHX
v3Vk6BfzzNYjP7fJkD9hFPmoUzCrNVDNCX3bVdTkmxjKGFiRfNPHYyZaiIvCfbRcefuSM5vi0Xbn
jYPGgwbqy54+ufrGuM8KgWMnveQyOasIx/qyERzDQUQ3GzEsYfaOdHrVwC7GTNPEEIr+oDwhWRvh
45MZaDQ2ZK7XLSeFpFmEXvbWviB7Gop5oy11AKH8NokbYKlJ2WBO5BwgXpBwGInkXhhHL1gXxm86
kn42bZ01vZaMKbwIv6CBMiGltBck/9gSoYAPb8AcsfF8vf+BZJoNyVyaOK2e1NVUB82jb2dvalmz
St5EfXSdVXfYe8dRCQFIsPzbe/f+lwTch959UYm/EwzdewAhUTXJA7hiSRbYaLXfrdjaKhxf/4Z5
1+kbqKZ84MfK0DstpEGwmjnMsz3Ho+ksaJgj/F+4LgQh2I76cccresAjJ2fcDbZfeZWBhtxQLkay
APOh5r9QxaqeIK0Ozlhrt6pHCiisDsMTvIyWRcNTbeEMLWjnvHMvP6YsYYGaEEWrM8nAmybSgUVk
o81sB0NDhIa1wpLLm5/49UtyE4rAHpg56D40qyujK5jm+lnyBrDRrjgliTnF1GFn7bbuLzkH7oQP
mjhhmSe9cqdcQXTB/H6jxhdiyPiY4c3oFGf+cV1aUrLa24O0MUgntc25d7pwOKGAJ8628ewurHkX
qHOy4QZReSAszM1SoQ5gQcdBbsVXp+1m5zxtE+DPEwzpYtGpbtTeMZUu1rvZFKDqlypYYCkN28UT
GAW/xcCiUX8aB1IvAg3fiVy0FBsNNfN2M/qLDcXh01pW7FLKKxojAhyJdj9lY/tGbDRNJSllfBLb
K4pnpMFejrjfp/LakYQmnKPSUYdyQQsbnyfFkDbxp3S1JpwDXVF6f726Xm5eIMrjRfMGsJMJduO4
eYdqaQMg6Lg1oxh4YEkBNSw0HBH9ocBi8vlguuoGNNeD2MtQ4Mz3KeOLncubgQV6nDQueQ4b2jrA
4WoJ0lM8B6DRUr8SglUVzqDxMlR90UTEJIuaqj2Zq3EA0qh1tSe963ASKbfa8eHa6mQe/xE6mJMC
u4APy3xEApRyuT7f8xHDmtCNHG7QjZ7G7AbMgIyCFAht6H8oxKRPswXqKQ2jSFusMnzdCF1T/ynV
HNCiP11m5tlch6rbk5LtcHLbx/0DOYWWOUNzGPIFzVLr1Qon91/x1BJrujoku/M6hArif5LKG5dp
ou1t9IGKqfUqWo0e5xAODGcjNruq71eLrHSh3SVYJEoCqTk283M2lezzmdFEqAW6d5JgHAn5McqT
RoqCYyFoIJXIM49R7wYsk8ohUk3RRsQpp+1lyai94BG64pJRRlztAL1DNtEFrn5rkoBUYAyneZuJ
wz5VEMSyGc8HjNSjRWgM8I7rPHaPKW2vQzMSWJUqLYw2Ol7GsgocZ0JSJBDNfUFUTlV3AAEIqsFk
lX2rEcbzUFMzvqOGzkg9hwxJv5nCvKDvrhBDjoWBrYhIUIadMpu2d1ocXWHdqjwr6eFZzWn6ClYE
sNqrUo1KCrIpfd1ft5RfUuwh+6xO5fBAHbfublyiXX19wpvOX9SZGS5DKwW7fh1qUFxoV9KaBv1n
3z5qJ/Qy8RmEGS1c8x9/pX0DCrwwHUrGHOgE96qE21I3+z8WF14E0GPEqhODJVqo4MZQU6DG9FsA
FMcActp2Iw6Zqo4crnFZ8RbnKNVJNY00iAsLb3iAWzFzF9Dzv7zuAwvneq2dnwfsNSTkv2OVN3po
UxReGD9AGvQmodgLPbJWJr6bOtWDSVVXT4UruNQbr3Oz+casdwA+VI3DSNTXvnFT4c3IFACdISYf
8x2y0HxMjpHmGLowBMUa+wu16spM0/EIu+ybvEke5FHq/OSPRIiIIbhoZvjgFFSHAiFp6yVgUbC/
DRTvkespOGIOaCV3D7BmrDK//9nmIK3u4X5e2H0A0rVeM9se3ia7695CGy/iGlB5GyLBLcvCWqDi
qrQSgjGFDgdDu8xlxgZP7A60Tb8pY325I65ymnnSEgjdVckLfg5sa5aCoP2mCEjXUzmGW9s3rx3z
GkhqG2/4MEMnBb/hfZg8iacqFbGCzaLaNj0opiCVNbcdNlOqkwhW2KZIhLnx/xfMBSLIwz3ZTD+F
AvSri6183zslGArLKjdok1onfv4uv5ezg4DpRpkv9imZ/8ISdI25fdotHCvEMAZblT/QS/9FyiSe
ZhHiMpawJ92kR/Fh7CPS6MOpnoFTo4bQn8r+5KpMioCwD8MSNsNMxycWi53sB1KWh9NyWiwe9uFd
SFnhr+ig372PWb4+aFxQ/p/6f6vYg5746/0HfMmf/SJReyeUnDLwBRk3jgg8soUu29qjQ7JxPkTC
6pe1dnAtJuAHDv0gWzUBARMqtOs06UPy9mgAODQNxDxHJ/hQGldx+yFdmsz60otKbOYMKCNIcugK
28SDa172rZz1FPOCWC6VsJMlPp/cw/hFh1bCFBcKk5RHWfmrgAnKOUbGbK/LM/KsiHVQ53c/iW8R
Fqdzl0nC9ODNzrnSZk0oyl6NwA2wrESfgpvyVP7w28YWF0C/U5Akhj1w+/ZFiWt2Ht8npgEIfGuy
TnsbjrDnKVx7/4xS0iUTi8Iv2cO7aismFplMbEFJ7S8MchWqhRe8tV0/Vrouv1neNyHlSaJZKQVN
i0DWGsDs7e7Yo9F6VR7EVokkoRGL7B9M2o9pz+9nvk/cFF/oMJZItuUbVwYef0hZ0vl8A1VeoqHC
Sym2+SlmFm0GUZBrePmIIgwNstdCwy123KnoJ0t6+BPmM0X20nel9jq8nWSFELBlRGgPlrTJeSFF
uQ+jVfelQXUimloa28sBiPGAUI6KSNF/Bd3EEIkyWSIxrS0lC4ohLuMORD9Xzi8p0izcAMjdnkGX
+6x8QP/tzK3Ogn66SzAjtaBynzWK9S0i0oJCfHsrTtEwSvlSsDRCnjgeClNVBg8MwlLDT3aHAAYf
STrySYF2tTOHiPgVhu1egtU42py+49OWZIofCjbGc1Tlm76N6dQVn8bMfvVqCXuxBc9ni4MZlq/O
QS7xDXdBnmvNqwROg3rhhQu/mjjXi9tCXEWWTLLHYfdJMiQQvXTei9O72as1w6RriMGoAe7ZoXFA
n27jPmtX2qas05yLxTobXOlEQP5APulmdmrC86ebjI+XiahGxfRKI2qxQUM2VS1z5di0bqbtAusf
7fsCkOYx9rsVYfo8claycJIfgP2UaRDQ/mJqA6mL99y1IrtrvLSR05YLaPbUCpaET23cDcVJ/Upb
LpR5aB9aqylMAuKRivtgykQktPPQrGSW69SglXKhxfxW1pkEuKJmA0J/8lZXXyZFrMAQ0y3Mu2as
1ArbKh6gXT4E1VVquaU5M9hJ3bNSa5ebyiIfLY8qz+ttRwow10VQ2aIeJAb5dV03JKqD9wC3/FZF
oDtstuiJ3YSPiGM2tWMUXDA/1v8T2fe4qXx6tSMckp9VDKmmhr+VEnLWs0yBZVx2F5nOSLq/60oe
23Fgs0e1dcmYUKUDpGaQ+g2SY5Nl0/DcG4qchVdVxr+rgKhDwMb3h1KLg2hPK/E9wScaKyA/oN/6
7S/aqf3UyE9ncZs9GDv2re3MauUebh/tQL3Enkt5Jxsakj4BlNktDv3cw1bzql4P1uk5vJREYq87
Xg4UfYXsMwZkjQt5tq1ikzrMxRxV7GqxZ++lnjh2m2s8I1kF4gvueH0+qNKKDIfieoS83m9Y5NnM
hXyWeRicaL+PDFE1WghHdAHL6xs3IK+QVHYRpIuPo4bD1w8IAhl8J+alEtnBc/GEhWB/Yy0XbpAQ
yvvYNu2TlgO8i5TBbyC29b0/Br7Mbd+zgYO//057FdAjzEcDE4m9OlKrR0OkZA49WumhW9AyHlSA
t1OV9na6hZLtEP9UqucchTAR5B5xlQWSUgmLJU5exihUY3GrcXCvjmsvSnaqHTrw/ebWm+Rr+FH6
oj34MAxJe/b8ze73T7eA3ajAM2v2rov7betp70qDKXKfUHBK2ftt5/ldsQxPs7vzF6fGjWvqgYtK
dB8mLZsbNGxNm7wY6EtBAcAlCv7y6sZ1YgWF4OsBdHEGrFD8mSgF03yD7BHS4fzartAlK83M3LsN
e+ndXrqShRi5qdY9kDHZjCGrvDtsL9zf6nkmDC3cRO19Mm8bjdUreTCIwXK8A3wR8045lho/Fg67
vb3Fne+Tk1qzdUmRjryZeWw8HNtegpldyNKk1Wqv4LPAHI2sn8QGemdlOWJ8F2McqipKhDVU4iSx
uFJ+sQE9EC2ns18Es+7RJKUPd2lUQ1yBnl9+m2Bq7SR1zj+Z29mlycNoaxdhFfdgjXxqTr+WyTyW
/kjBhgGDHPaSLHl+BH/8bqNBQfDWaxGrRaWR/F6FFkxZ3gale5llrl7WEEeuAwC2D6jKCQ45GYoz
QIURqxpeF/+yfxySjL/S8jzVd5zVwZ1aqgev/10b3Px9OUoPNfIX9oq5MCAD7QLyPXyi09K4Wdbl
HDanNJea61br+wWlIHjWFRPX3oRhwihmvbov0zCpRou2S2gZFzrv3FuPWiM2+4nvxqdplXXHoBIt
3BJb+sGOrjyGxbEYE/vffFJEEKcofqzODRsFo0xYUxNhD8PIerejb28uRMT8TjvT45p4FX7Ik9CF
Or2qAXbGoCah4DlUpAkn7AYpJKqeP8RwZjfx6HsvFAn4bmKiAtjSWX2W9T0Al7Hc/Cd5AqfU0/xF
l1BPgHjlmtoP22aWYfShL0T3twQHZz7HJp2dEK8PdeulyTy0OB4SOjsbetlfVaWng0IcimJq+IBb
b7MVQdNTHZIs9s+Hkz2WLKcdPuElyAMSTRMndRnsBwLWhoqR1fNqwJcoLjYLr9Ub5Q1gp3lykepy
KVqa2RhrVVixGQNhWNXlQ4eHmThTOkGMnYumRF7CqIj3r44oyKOpdz3VIJsGrmiqSG1g3vPdNSJS
FORlGx+7Z53+GodKpQ7o5CrN4cQX2BQkNdshuoQCC3JI6jRQFSD5umCEwqSHCT5Lv2/Y0JwwgqcK
VQvW9hYqpeWu7/oTOo/r54mV7YnQvBaLlCvemBCdjX3yeBeW//jaSnv7FcfVQ2vvHq6xqfa0w52h
RtEz/vLEkKHUjsWp9ZElggVijlpET1OOuES4hThWUDqZF+ww7GozE+b5HhIVTIi4Tiy5Cy3pJKOG
/1JhlXqBaR2X3AfoRBDUMQZ8cZJf5sO41IGkRM1IFhLmoZRj5NjBC8GABgeZH8DkRV3WQg5ouhjR
YXTpf41Ur7VflqXjVX784/kP/KYsuKh7EYMLbbd/qm26wguAcG9TCX1EtmzZEEqzC2TT1GSV8wZm
NtQIFYu0TaDW89JYb0QM9JQh065qXygfsF7HRVSO3AvDExyAMLv54cqPj+5Ru7rtM0/Tj3eJ9NnD
lIxZzeA3I6GXoF9uzHv9Cuq6bYXSDFjhozEB08HAkGquM5ID+itywz8V0k4PPhuErIdzzhCvmX/v
qYYff5PCP4/g/pu7A6LURE7/op8Hx8l2Wud8ZJGlufH98UMTZI0W+VpgsjASXnRodcSpm+ejPX26
QsFm9JmvFuGkbMQbOi26ZJbDoV0v6o/btVjITOlasnjTOkbJDNojwV4LKjm4a/OAzgGopYICajT2
57Jf4PZJLhOqbet2AbSTFdVNkJmNa2ECXo3SUkAgY91LWWwmhXhx0ORyz9m2Jciw/SzL33c4NSbj
0hw44MKGV0VXAM3C+6yd9+gP+UXsKFb8qwjViDvQ7Zd1QoNaf1zdDNiuDtStQxz3DwGn5E0U1peR
95G4DdVy2o9LiVLvX3DBypwSZkLlbv4vCciNVJwWTg9Xbk70FyXOwg80v9hc1jabjZIdeGCuMw3Z
RiW7KPeS6tYbowL9LT7RPikYe/XiIlAAhdrowTP0NvvDpoA1RwWxXn/ofeuJ3pR/MgiDbx23vwQG
80C0Va4b/R5LtmKVu9YNz7Ww9/bs7QE0cPQ7JosIliEwjzV8GIr3kl/5IeU1Btxv5Htmyb8EIG9X
+ZYkMrNEkVJU6w5Eo+70jwgiT13uqsFPDJBsnn8GUAWa+ZOUXu6zqlJk8wdkI76lJjbrp8BdLsh1
Eb/udZ34ch1WaO5QPjDZcHT1PE52mXDezpmMz5JufcVoQxHvXRs0X7Zy9ZASCpvnjB3xAL8nXilF
ZMWOfRVA8Kf9gsooHpK0gF0GUKLt39Yyk9nS7s47u/0vJjwp+R+gt0lTbCXkjMejSnC4LL9Vy86E
BYY56aBklMb8CZEG9Orcrsi7bPmZ8GpjR5pJ1Ty+6ph5lMSmDA2MZBR9h4sRh/gLiiASleVe35Fd
wmWQ9qwdaUu0uE/+k7WqdjNbKC7VupQfM62kKhmYJeqxujUgcXMgrGMDHzxMdCxRF6m72IYI0nlw
k1bUfQ1Z8NyjB8Il6A88LlHBZEiXPfdsN9A/TwlvrLo1AfipPcMJ3yO4VfWYncfy2CHZ+8aTQEvA
tsrjVKMXya7UeZVqttv8gwu5de25/nBpcaS4SBFvtNgLgM4/WkVcfiX1au7W7oiJnEsJ1mM/fFqj
OXPHNPrR60V8PBGLDA+J2yTWZfwEhH16mYLzlmy3TDXO78+b8spLCYR3Osk+MPsG3vBETe2WkTIu
OcdpLRETXVPEfTAcIBRCI84WSenVD/+3CGpyNlvLcyap1Q9ZC3sI42uLIXP1n+F2UwbvAPX3ID4h
HUk+fi+Adz7wF1vmx/aC5ZfgzXTf3JyLbxABPISECRwazRK7ExSBWUUi+kUMY92e1R6NcvdyIh7A
O7AsuTrn9nPomG/0d6qnxxLnw7H3ST8GL4UzLw2nnu9SgY4zJBWrOy9cutXOAELCNFHBK7uF8ljD
Vq+AnFhZz2evpwnWl+vGi1QbZJqM9MWv51uvx9dwKH0sKJNaX4AgFABQpRIsi6NQI675YTaKXIqy
3FX68njXi16/uparEw672S/pCzgz6PjG9KPmjSbYlyedKbF5IVKFIdilcccKzbZ582b2ShluA/Sl
oOXYFCA44g8rqiwq9AF4mjswx4cNcylwYylbF1iP1dmrnRyEGeROg6l6mVdAkwkRl0SXMA7xdG3d
SeyXLRaJILscUolzojAKuO5I4TnjxeHMVaqA19gRIZRpUiJin5maH/xVc0C+pPPhxo4z10QZXCvr
TnYftEMACSKaDARlmr8unCbMcILI4iQlmemP//otudwN0knKusOTLre3LujVsURMYdu/+wA3/JZl
HmvNJvVb4hsj9ol1l7rP35izG90+ZLhN+xVcqERSJglmfYnQBFVDfR9Cjf14tMjrYDfqkWhz4XjB
QefSXl4kWuWAZOWWITsexhhAVyETy5dXILUs3g48LJaRNLwE12oHZSF+KeVhmgpDXfEnDFcLYvk2
VYSKZ7YJDzMpmUHMYJ8HRpYbYC8FbNZnBGY3apwhAf31vqPQyKqKwzIoZVGhWEDSwWUc+8761O8v
Sc+ZKmlsuqb3aFywbnKu7sdK+01zq/FsME/AJUyu0HSjGYO9AGSqEzbTFkl+9MToxOMRseJ6daru
en/nnBVdn60+z3l/S36i2o4xE7EUkKfzJUp1p3qcyqdR0nXUT4SowSdj4fhOIu2IzPrLtVCElVqk
OqOqw4zD6ziNFIANWSTP9tcoxeJZ9ZOCsSwydrB71uzO1avl1KxoxOa0nYn+6l4Fq5+TY5g5vhP0
6dLHdQAhk+kViZbjgBI2+Z6fEEsLcPav1pAp8loaaN16pwNX9043Q7dkuip6uH2vnGgZDYha04hz
XHrKc48dLDk3Pl33GTbsgv0VIhbAAmpT/WMs1mpJ709c0yRh47b0vWdAtLIoVA9FhSEOIyzsrYBk
C1acnTbwo0nw77NvSA3P7nrVl3cANoCPtQwCw/CmyyFAL9MN6qGFv34aDZHV7wRjfVXb1smSQsn+
zvovxQJntis18NKYuj7DMrt8X/H/TQ/9R7/DA4idbPwuXyveQeIWCsthQVKT9pb4KEwOYd89WNnm
WaE3y+ca+wWza51FYR0g07t7+jHVU6LWZJYxR2LJf5pvSAyQ5peYRhOlBYhc6pEY0qBzQ20CiUx8
9hINyTk/nv350ONQTKKw8uxIlsE9ezNjaAkPFsHoU4Hwd0mp2rUQUgvr6qfJGtMmMJyBGytuVovz
9zyRg4Ap5saXB5n1O/+J/CE/4SEiZ96EhrmCbwdWSRtgO3Rygd7EmAA4vjLq0WUOGf5KmHCQGc/x
KZVgW2NX8DUml45inYe5Zk/Soh7H0aw9d903ewy5vSNPEfgvnreDokgcR/y3bcu+AIhDoghnL9DN
+UPD86EnpaAON4YWwrTgewcSprL2jo49U3Lwjzox909n95DKfc3n0u8/l+OnWrzknIkhR7SSn6Mo
KSjC5H3Kgq0MgeAF/aukhnXaF5A/wkYzjU/EGDHOa0tU7ifPxXM6W7OCtDrVzCfOBAGAt/Ov4lnd
48J9vPnupXUbgm1NH1Q8tgv0MBZO0EeTaJdjSjn/5hMhcZZc5W4Nz2AixPHNzHyY9E4mbba7ePpB
XtYWVl0mCl2z0GROehGq1IOYujj8peqEWmaf6CEBZq+eQdFjcBjn3OQvaY/T3NKaM6IYdUXTZiEl
pQAcQHUEzn6aMm0WA7tGe8awZJwKzqCEkjjo4U6sR1fN2Q4RbQv06cOf1m2CUy1zlnA6g0p2yCJw
ssN7AsKCk0XqS5jRLn8+JO//PjQ0fP4E86GBB4+UZx3cdmJhRjjyViV4vRvy5fd37snBBRfeQ7t4
CSndbybNOS1p4PMrejTI9JSALUJvPadMksTg/B5wFmSFE1e/JtmOv2SZRkw/vfSjCxxBPXtQeH2m
w1LDAIL3R56VQAMme5Rb6PX6G2wBqQ4ga0VGLQ3Y+NP+48O4c/KCHjXwlAg6b4NsiYHKNTKLwjSr
7Cwzf9cWHCAgJRKUf6LczPuJE2/PAtQWC8OZHUGnvteLaByXX4cH245GiQw5Ab1Ps/u8ADl0HCOM
lT/jvnDiKTigGK4+cm2p/gKvI0VlzIq7FoYCGBVheZps2gIIDYNiTKxP/xbrbQXLH9+JomIeeNHx
M9pwtqRLDm3Lltr5ZJoJ/CvssJjOGJXe5W6T70Nzz6ExsI+kK5g//Qqmgk5a6GWAIO50IBY8n+XW
/CLwEzoA7nKjgm+jHRUhf6O1+ArAHBMKheBt+hAIIAsDLvg27UVjeys2xU/rvvM5ESUcrBDKKlay
omyUA7hWRCebajPg7B2OAaFgzCeToifczB/dQFRsdSL9VDUtX32QewEAX0zBX1tO2v7rLl/PiblZ
VlneLZ4iAw58Al2NgnaYlFJJt6xewFF4mfAAB2bwlUS6cUf7fwoM+p2pcYe9EAglkHh87g83RUYU
h75tDWSy/TxrRL4XwqGwGoeXGyYCfYNo9bC4SZYkruHj3ljlCSkYdqqfM6mbNHjpIckSCVT4Vqad
jjAUiVVcmsps6+MTHCi2ZUM5WFnGQkAH/NTBOJkq1TWxgSG1fDYFMEBBb7G0jC0Wv3UrxVUvujTm
QsQG4kROTy5HtJCOQVeU5OcszgADdhRRw58TMHZoxXcCQvho1FtwWjefH+TLTpFR2RmpnKdQDcHb
6Oyolb+7Y/BVgUoC7rCWp2lvb5PK4DMdngTd11dZeX+SWaMiAVPuVHTjq9nfjrwiFfkDNSd70P2s
gsPY12MBdtvxItSw9TEgzdzQJll9jpDsknnJtc4BWrFnpAQmjAvzJLtt4iwy+3MXNNcXH4nBAnFP
O97BU2QG6gCkuDNDI5gBPiWBfDpdqC8POhWB9aSNbkRlse7y+ILP/62uM88uitJXUpqhZOloggpT
0BN0CIDKL4SGA+JO7FD7haknfsm9sCffpne1CFmhbAnbUeT8h9bGobvREsGGHdlaqNCSprGxuAnF
LOXO+5r2B6x6AGNX/bZ2p+El7ET3vKPHNQ9/BXjkFJp9B4r4n5youdnISZC8PE4DZ0u98I4bGc+x
5pHHri9/Q5n1TOr8/N5pGz1ATYH4BFMMJJADtxmAESAvRt32tccJ4w4TR8PzGU9I0QLhlnRypcl+
HSSRZc1sAU5XoJMKnboyzT0g+era109RdMbm7+VX5NcdKFrz5FTmqDBUlqeftoYx5VpT7TTPdBkr
Fnx5rMA+rMvoyvsgl6XSaupCj7a9EeKa1XrIhrsfo1x6fsGOH75unPi/PA6IWEvqJ5QNUZTsrr2O
lXxjekr2qQI6rO0WKISn7PG2om68qNeTqZoBy8qwMo6/CvWrunabGzjRf6NpYvqv+baoNM7+xa4B
BMPwE9KrjC18ADRR01s7Kf0GjGk+rHr9uI0UNvj86KbmhsD5k/SYfh8hjVS4S5FeHGbmdEDkEZTk
R0rrFNVfy1vJbhlIMNyK9wLMuF528WOtjfrqsgCweKNuE11911brWp9e4j7Gjdy77vCIPOIlA5O0
vYsyncJuXSsFSMDPAKWNdlIqf4XOG2S4zIx+1Z25B+w1Wb8FqAZkwxkmDa7S5a8JAyuLV18XpLol
Rz0QQ4Zd1Ui1Pgb0NcK6qPEcRC9qFjsLABhi/sig38wZXxUgGVq1dm++r9mbr1Qj40TrwBeu7Dwr
vILoBLCODZLsNGCCpkal4bIkTIMoyeINZq9gsiAZTeWstyOsPfCLa4fB7GBSO+eHgl9f7bJc7De9
wum0F4DIt5+QetT7JzRMqv43qAqhDtivO0+EH1qHt43ydTW/BBh72lEv8jpv//I/M+QfzuCa93QC
XP9c3e3XQXWoG3drkqPFInu4KsmOvrbac3CWjnVaUl0gjff51Vk1we37+2ef+0Q1Hzh4H4bDo9+5
CWdygu1fngRUMNtEfHiGfMfSHo47pMD0euchF1E54M3D8ZGVk+aHByuTH0po8DeugVLStS+GfIb5
7f9n61L9AsBmSfI+myy8cPhXvhdqUQSB97JZhW2EBHBK1jnZkL94sRpApcmxk6jRXDeQgX4l9sBH
uh/WKbqAY5nSvw9xI+P+eYGMjfY6U5eYPBuXr9PmXmuILU+jXKr99dEmcU1YODUevO6JK5i4lCu4
9rATYnZtapfn56X4EG9pEpWReQ8qxAP1p7SOlz+oJWI+WwBpVeCHoqWQUK6j6c0O0nhKNIRW4Dqx
ygmbOyEICJbMEl+kbShVw84e92sbLmV7mp8PlTU6qtqSMDe4lxeTJ0k1c+CFu6auQbpwyg6Z9soy
VanC8XJZNAPTR784c1CKRPEdv223XbanhKjid66l/70fVTkgdJp6TEZdO5OHfw7mVxISLO4SBLBF
pW3RtpzGzedE2BmjyjwIIzG0TDYSaa9x3wvEpQ/kRKqLrFSvaa1ceHCFFuo11eKTo2ikktCZ0VKU
23p0ih0elc/qnMr532aYGJFmF9OUK4Gc4OrL0o1Cu9rI0oIhLiQbM/DMxXiUxA03zEN95Z9HMx9b
FIVslIJicP7d9kxD/MfDHePJzOKhU/uhU63vIkaAXImSokHXhwtw/6PDAnH+EsQLhVZlpC23/VIF
DPcDpAn2hlCa2/vnWAA+XhrHtE5817UNDzrQVWEd8WTC082gElQJ30C/mRiYO01YBEGK6BMB4bP6
k01xMiBMqSAlucbAhzUFMxF3CI+h3O+5zHaFmKhar9wq+RhM+M5FU4EnpT8LWt+0B+Hw7zrm9k0v
k2+SObP1IhTcqCWqP30lv/z584PmhzXledmkn5x7vjRvJ6MQ1okE/TZg26yUWW5IJrDq7SzFsgt7
Hjfti4X6rLcJkvGNPkjiCqMz0Obh4TOIAAMtlC3IuZsMUIPaHAHWRL34YS15jlOUmmWWuHxMbX1x
BOcExEr8tTQBrwr3NFSe9pDU8412ddXvc2NmqLMPVwhPuX/ZvzUoe4N0LOidvErVCyWPAZq4G28X
MMy0HYlMSUQ0Nci2NzJoBLcNsN++lWMpKs/o5t2J8Vf7Jz9f76VUiKtWxtp7En+WVRJ9ZCQo4tIW
gc9ZnIOjouwLhCybFWzl9v7gEB6qpHHTofYGn6pSddTH6z8BBQCESXTH+4t6oP4Qz/WAXF65dXTZ
GVfrDPVRmCGQfw6An7PmzQ8xU0RN1jjjegbPR+xIJamRdJc8DW6JTlSQMu/lsiXZHMoTzXK8GdwK
kQ6ZNQhDvNVNMExZZ2kiQ6GO95N8vO3Dy8+K21GKDeN2gS+4E4VJoXcnOjXBDzJsyFnc4TlBg3xR
NipSbW49DnZGQIVOzACxMDa21AwGOqszyRx3i+b0Iw+iVwZVXesNjNRm/zOEyJrq/DFiMGY8hhtU
74+g4m8hD5/ImBNA9NcN59BxJW+42PBMys6CQwSyS9Qur+SR/gHnH8eA09ah9xVFCzAeWpVWy2Wm
f68ITtE6VM+yMwfFIdqq9wkBI8R+u7kjbHFoyeW+ybFUbiJPX6SG3EVxZqJvygJpE+Elw7xLlCK2
cu90Irn2db47CREXItQZWpIDi2aUKAREAUeghyc69d5MIzuwUSWqkV8SoCowjeTREJSMFsSdVHCt
l5EFiHn7vfSzAIIKQ/xLFUBlEblbrwSG7tv9te0rC2DqnrSxKH6arhezk/Dhps1y2Q1+SzW9Auy5
xp0FNCbnY5iyR2czG2kSs+ji73DV1qZBLDD/um2BO9afckr+TGqRLSSlFKimtOWkJfQojTa7ov8F
7g8gbGXMFWKCTwJrhxyjYqEdfboyWfHqm6kA7S6H8zMhZdb77Vtkx583a/hUDo9gP9l88NRYafLI
GAJbajZMtWHIaTqn8MFmHLPp1sXqn8eghDkmjst6JdZ2lBx3hnR80FDR1QiOsG8iuHDQ/vaS5BKM
JDBJR2CV8m3xmS3aS0pO/JQUV9xcKVktJErbRClwBrzuZDMHEPuwHkxyHpwyfRJQ6EiL+qi11pbu
JkMz4RRJNpKzZ38xAExW9uGzVND5cvgsBjb9H4nZtWjBD4gsUq79oSsxBMW8md/A4XTs9BjCWG9s
DGyujm8jvgYhDuPys7cRf1q31L1n1uC/KLdO8CjzMY+XBqj/ZCKuKIG9fAP4fqXqIYojxatk4T5s
zSeAFAJ5Vq0U8NbEptrcEDRic+ntXBpFlIp8m6+M/PaTHI7SINVta49FkrIZxhyOwuTAtK7n9ZwQ
G8KIrCwS8VoLnr5OIiawW9SjokzjIieF5P8uawecPe0JmKtLpLn4bwE6+4JUnga2F4QPb5OSg8xB
nPt/Yfln7mSYacztkBYYB150vy4K7VREobSMyqJZoc/rky39ijxiKVUTdsVmEYK+Wh5xtBZreSMA
dv02sAFbBp7Q+haGikTZySAp9n6YIOc4Jtpn/1ft5fGbWV3CAHve66K5Ol/buF0JDaBvJaKtRzQ3
Psq2GOhlNzoRBqLIMxzSpnjI43j2pDsLKhg+3cKT8IBL1rFXHi9da1ZdOP5flmL4gp9FAAusxAhj
iJ/22Dp6ncKi0xydxb35C9qZy4CdC1BWokDkbCa8M1gD8prBdIlK4tWlW/LB9QPcMlvfzG2Vgpja
6K4x6wi/RNuSNi9Gua/Lhwgo4iKXmoXIVP0KWot9ikQbCDgeYA9ntjoegPKT+/nWZSR8zTzAvsBF
w2ULxBKGGqLWvEYlHaS3cPF/qWBGO6c0TnIunin1FtzP3kxgd9eI9P3uArkgHamsIX3od2iQ/0Np
i6+bKLZUdE22vdIEW01JroV9/Ra0H9ojW9cYk3jWNSbBuIJ8ipXsYvBu+Ios8+OTG1eHm8+AhF+F
3mQ8a3SBJbCPBY7BTVLKVtkFiLZCLuScPjck7njSOU7ttRcWAvIW7lSNSh+9FhOqdfzYusgAduA3
gafvLSY2YA8pbhoFe5Z1UF41V4ZLnTiZlsFqmNxDOQHUWL3vBIuhkxuwqUEuTd7Gup4bNMeedQxu
6Tq1AGsGxzBW1t2z+BTfRqa7710oLtnG5x+Nt/R5PSrQk1FCKwtmpzyC4fT+mWb/YkTJtMSv8Bky
F4V3HnsK06197HMJ2+3Gx/A9ZJT88U4dm0g4CvPPA/A8I/fn7IdPK4F3NCXATfxXCUs4qBhUuYU+
dHAi5xD2jWvOKUQGLHCGWA5Q3gfhzKdw94CqBNgjGbrCH52yCXo+iy3/9/4JhqA854jSM50pQxt5
QSpZmEtGHA4iIJnadTQ30jDYCfy4er6uHDvbneypqSydEk4m/ywUImZ0IHhNvdbMXkJ6TqcDFomB
qP+4U3OqVoJBjcUamvIZah60qTTfrFexvKToTppPwEYESi6vBqM1abUb0UAo3Rk3ApstjvsFFYaK
iD1kAR4ZpxF+hww9cD0meQOJcxGQYfx1KTV2HrBT1gADuZelaqIAUMbWdqHUFh10//S5wdwKpjdv
NfxKPhberBCucZqEzG8/g+A0SnkT3+jyhZs/R+ZiXn7zPxFN8qERRPP502cY6xq+xUDZVB5ZiSUH
0BNgajCxbEqD4EsipSVCmKiWuAK1Yt7vaxruRh0rBQ5+W/xSa3J6UOColiltNkn6WoiNIC4wZOW8
aZsogYa5E/DPkDjDgKuJOjy8RtuuJae3guZQE5mzscg7e8Ly457uU2gaZSEnykj4q1nR0VwM6gD+
NRU2o9v2hevuoHLG+l27EW+9iwBU9275f97bNB2KmRJb8Phatq0Kpr8VuI+TfSNisKJlIrb2t+DN
qMoUqaYi/Rpp2b85DynaujMmw/7c8YKhvQQTZQiRboTRu8su8i9Ay5WdM6vAK3Wj60yTqv8MdgAn
7dHt3pzgjgLSwAFDPoRP7l67bOoNOliwjHha2mbn0FGg/qVEaLXrZ81eMPqJs79Dg5w2LZ2LEELe
sLVghO5Ef1hfzoA3OWAMh95Kcu5bsYcA2veYAmDTytnn0CSU+MHBli80QIhcG13CJC8t67NncBzx
0LuZ1V6cHnOHDpQf79y//rfi6q32YJrHhhAnXfv+xvajvtGDImSH9KaLqLruoecaGz2kEQ9aD22l
mQWKL9iaJfYWifRS8zt8FZuaK7MkzNUBvKMYz6JzcW3NwBvyTviFGU4wSvAA19yUImYLAp6E4CXk
1CLKlZXSNiK6/m2pf5V1AvUiQS+I05qVVhfF/9rU+HA1EShBa93HQToQSkWiVPPMSLaY2il3gHVS
pFMnAb/t3yVXN2LFrT4mIs9p5Oy1a5MUzkyUS5a/bvRJIU7RYnrJRaMW+dD/yZ2YU+9aKq2JNbFx
8ZgaC6j9usm/znprWl58AnuY3QMC8tLzlYLpOLUN5SJp8oK7mDGRXAz5EJF0tAo6/mb0vSZCkq83
76qVBCWkIWsS67911yXLL5DyR1tvwo5BkshC30PJ+JqABfd7ip6AWzttx73XLtSNWGdHmDC/y1X5
1rGkawOgN2MiJiR64KTtwB7H9uSW9xEOp6y8s0anyRRWcsq0yIBgLShqJSh8F5ADDkgAlKnDMOkx
Ct7oP+ydqeLrKSfwmBC8UYmVn4tjIzZQZg/Qbxq+HOUBvuRit2rFGuesqEChyLHKl0nv0hcGF79h
uE+8TS6OUtF8DWojobmPLH2cG3RA6XFdJp+2QfGklry3cBJ1o0V32wg6lfX4QFBddmxv3kQ9j8/V
03wF0pTcx7kuufFNKg7P0OrbuCZWtoGG0uUJjGGM6JrGfqzphmiblf/eaKFk5f/0YQGV3kauVtls
etDxKrndEGIoDJsIGADBwg6/PnIKYowNl+wAarVFT/2yQrvmrFPzUVklX/QxLXwrD1/clnyQxzob
ZJi/0Gph7RYZpHd7G52y7h3CT8V6zEB+dX967iwn5p6ew/e6NhMnYmDKon7pYAMrNNO4jlEMQs2/
zmPxAgJDGoWcxfcFveYoiNLT35DetuQjJRC5FRDq/2ZY0oQ4Ofx+6PjVKTgCERkVUV7FbELuEV31
HdvaKCCI4T6fjjNVswRGdQBpQOAWEvBz/zyVxa4nqBpqz2WkDKq4ciahnSTEInkT/IZUqk1520HE
Cxy+1N8eHFP5bY+EcDeVLKIM0igfeBK0iV4pOwR+GPJRujtTqnF9Gdxs+kK9ZjA4sVKjGoW1+aqA
FMY/g7/WUB5G+VabrKX6/UHGrAu6FlPZXNJCA14+s3J5L1M29CoG4gjH8Sxvec3ZB0Wa5lvmRCht
w+wlktapqyTsdoyzJw5nhRrPhOfBNa9HNmhRZ+kntfuSxNHVhLvN/VlQK3RtrqHBaIWYPJ/fRT/m
0rmtwMD8/ZDK5jBda/vdQaOJ5Ibp7ymKjIq7BdYjDlBKxxOMU80umzPYQQ4riP2c5Fiwqe74nVD7
D0Mxs/nuA8xWI2/qHLhngJV7QPm2bgWtDcGljRHE5+c3KYI04PUayLolMCDLUHMYxSev6uhY/vAq
ql9R3fPGwgdIY919FkSFTsES7rv0h3ZKHGtOkloDwBWcycBVwB8WPoqQGquCdx539HYDxctgK2EC
73cLkUFhJysZeHmkvR1+RGmYtc5qg18Loxo/F6cWJ+w2hOOO5FsLX506JA5ExyTrKrtNbZbSqixT
gEpf4MfP9GTZyXbGj/gm3P8a7LMR3YYXlkEWNsusZ2u8yxymE5h1x5P6fNyoJAoJQ+YcnGECIuCE
g/mF6DQAyc9339j6ZiHvvfv3wM8ofEacE6JXJ7gy6RlAxWbA3XRfYp2W0Wu2ZF7fTjsHO6xASaYp
K2u+56NLmEArnIRUoDVFFZWjOz3g1m18S82DA+A0zDQzW3MT9WDPv5xcLvzFpEgX+3j3aF/YMrLK
VFhM5At2jivbnbrx0wNooEage7/ke7qQuHD6CmXVOqlDmYdtOs2uJ41+iaLdS3IV5hZ/Y/S/ycky
+qMNKBPZ6/XP6KbkWU4ixtZjqR1jDr075RKt5LfCcyi5DJ9CGyJji1iab2n+Q/D9q0vYb61jEK9g
MS+Ir2FqwQZD32KiAxdfJYGdmTPVc0C1JFNI6t7gF9khvefHcmK4MIeQii+smiIt4NBquAOs11y7
/D+RPHrqTweAdblbXT6HJSXFtLrMAkQbQ6qEzbMf38FdMbmeKwCc0zBxS5dlBcq9Ww3WYfeE6isC
qY3T6uk9Nrjg6aphQMMPp2+xYNVb6ASa/r1TRp68cE24JApmagwCg96nLbGjBgFwZD4H79uZA6al
gXBKoTiBLE08TFsdOkGRXyYlMiiH/DUaRI0q9JDWhlqWpoOFxTQ5f84RNoIk0sjlQV4AGggMW+X/
+FChVSSEValX0ZqWnLJkgczwizFFUMm5QvbGkVaizowbTEJ9VBq3IkHHfI6a+Us6yDLHklPI73Of
AbiSkg/drJg25jvE8K+QWuXEb7poZfbdOVEtKvqixcjoa6k2zE28ee23Ypx82U1w83FuuXVZplLc
mq0eF+Oh68bFht0HnF3vxUvZJ4R39pd6ACXnB0K6RK/XgJ3f/0aTJFqaNILTYGM5CDCDFLmtNdTV
3jjqm78a63pAfduJ5twXZzdVyFNGYV8WmVsa28EAINiWy3mGhctslOZ3xkirQABrJuPHjLUH3u5A
1F7mJeOKQ0Rv1qU1D44TrlklFRznB2LYIK6rUipIpKp4QLjm+3rIDX8ydGG/UeqWBpXVLmEDGKua
IpPADWeOh/EKW5zXt/Mn+bDY9xNc1tdGmPXAYetyRivOdP76w/8I7IDLK7gL1I50xeEoR1ADtxzc
os3R8PDJfWaiemCi02AEPlfzozO7OzcCvWubYFkjnvtlcVBsNCnu520SGNgEtsxyilXlz5Aby7sC
npW3K+rCqNsO7PouDFE03k8NmlHwlACbCAHSxMX/9pgtgmeXEVnHO2qRJbxF5wuphk6HTUr5Q0gD
jTUHmEudSA7oD86nbkPgGEnwc4WilrLVl5b5CUKXqJfHhpGNJLpps3NA29GUFTEFlK/OCTsRKjpR
QEbsdB7qfYmLrhTKq5t+m1NIGvwmtMTFr9E4MgSWcIBe4XGpEboepYlN7eSFjysb7B5KTN8TYww6
aXqsIFD4oL/r1XBOE7SJ+SqyvaiZY8ISAiWDzcmtUuaiJLkgluhwncNZV+5TQtNJeA//fLdHSAtH
Ket6lVk3Mya/hOlycoBNAbwUD631BCgyzVd6wQ4qxPBN/d7nq3FVfIb//38LbkWYOIDDtYWXtFta
7PPe/2VskKEgQC9UeBC+DWuL2AyqAcNDuTklywePfwPmrNb7wI7bK8ZUCTrU3j4HTnenPqIW7emU
NgPOsRUh6BFcWr7GMdP0BaQ4LiXkglnc9+Fg5zn8EGMmlHPDkZEhUPVwWf6JOfJbxVmkap8Fxk4m
3vFaEcbvuaRwpXQjQGDfEVt8/LDNu2AdGAPvIadVHxdzOwLKb1tkxtqI86ibKTNJiHWa/GiDv/aV
ARxClS0mJbQOU4kYE1nkRMUFkm33PpR1z1SozswfYHGsq4H5fbG9HWgkExUR6ECXWLwSfH78ZwXz
5hnv/wiYebgB5VXXy+CxPzuA2KUghtdJbga2Q4a/kpQjGR4lOEoWcxmkxRI4mJJ7R1fj5wWdn5sZ
uKy5dLAOgx3uOD8p/uRGP0LNl0f9/JWzTogmIrH7H4M5YWlEd15pfueSp7ZAoFXIJJtc4eDSFgqL
MIxRHTT7aS/rFurxlycG1wa8Wic1sScDHCMF44KJFeM4/+ClxbDcsPSPVfZ1GXuYd0m4IeyxhG87
dQpQT87EcIqLV1IIjYO1NsXhwleqy0Bb4jtaRgemQq8XcuVzlPcN1w8atXK1hyQq7/K7w5lyOuM+
CsG9Rj/S2It7pLRVJPdBXTK7V+ip9BUBfkJ4E/xcX7hsEuD5vTh6xc+pMMlWMn0KuFj4rbrvYcen
r944q8Z5nTlBITjwF718SI/TMoH/njESsznND8SoUW8jkkVlhSuQr9nyTw3uw1+qwq/gULNXTd29
QWVUy3sa3cmfK9kz2s+Py4BFWcqRZq8AkhDioSeNnbB93wMTnmqYCMsAtz3rd5muB1buwaGJ4hwf
YNMi8mQs8mP1lqVDKOoa0Lgs5MoOEXiabc560K2RZPJHOMwgLJt9wMde0tbG/oHuBKIrZwwbujMN
HS+4NRzJP5n0psMG4HbyIwR5h64J2o8znk6hPCpo+6fUnds3AZPa+dVHD3hQgJPQ5Dya9TjhQA63
Rm5FpGrxi2WKHpGvUrDMO8M8wNSk4QxmAwwyps+pa1vOuzXzTRr17lT1Zgm4EC5fpEMpwOTOSdrf
Z8eLuCUhTQUVf2l7TU1LBYSAVn8YW69dZMF6/mZJSB58Lu5UPqXHDuCPY4WwuQywOEyICt3stzBo
uKxcw0cHvWZqBwGxEpPBOseTzloHVUg0OGyG8BsuKrrEwz7Bov9qoHY3fYb2fZeFplizSVixbIvy
bNERHHNPn0T6aY5HqCvPSr6t6tXjJ8NdCVKkERp6ANgsfIEorH83+RhEU+Mq9mKMoHo3YjM0/Ha0
D9M6+KaN37Y7djuLpeTthfnMv2r451KXIY/CY8R62dbrpiY6QxshYvXEHT8eLt8pGlrlfN80EiWG
MgU1WdDgpWXrdvO9q983kYKEeQQyRovClrsuCehSkmwRuaCGgraZpPWQs6BppTmpVsQf4ptMG/YU
ghM3lJzG4f44PXa9xQWyK7ZvjhkS7frg2x0BopZYHla/cikSmIhH2JIrvzfRDgFU2NUXqfx2Ad7V
U4OlswHA+7AYvUPCIcS/X4IXKk6k1u6t9qo0h7ojTibAbT/oq9dPiGbhF2s4rE5RlHDld6SKsuy9
xkQAGNQwNOGzovx6du6LuQkAc2AzFwlHYXMVqo4Wp5gjTQLCjQUNh/9aQMyQWCNse63xVY9MwUPp
gtLZqibe7snrTOualuReSa1XgfnUimw+WFY/ciuakORhfT8IQjX25AryiaSKiV+OBi34tsEi9p3+
tDs/r5W1wShRx5nu6+oGx2o2kwRMnlFyQI0wEJSekkK2SmWXLwoY/GtUXNNdYa/ChM38wnpBQht5
t8P+FLCuAmauqDTgzZoG39DB0/LjTzn/RwcXK0V7hqoovO3zDgtTMRkwuzI6gVckcs7EFuB0LKkB
VlT/0JaRzEwWLpn9YcuVSCTnYapRBpr6w2tzAn048adedIAmRmRteg6uL3zk9DrDYl0Bay/kQHQm
48ipZwAAlVxToyerJ/y4FnUW1xDr220lsadftVKzhV6rKfJmxHtQuBD56zrgoTLgAjdMtw/xwupA
O3VX9EfDvLDvn1UJ/yBgGWsGp5n9NZiOHuvSJqlmnNL1Nisd/t2ygYXsQ6AKQKNCoaAm31Zp1zlJ
7nLdUJGkJZFRNjMn7CULSr1WIJGmIekykvJSsX/w/9m5bzGvOiTGKle2RiNPseLcjLrvvsjACWA3
PeZJE44QwDHrnegEwWKKD7hoI5lHZgSrc+r5lq7ty7HppbkK5q9wPwu9SNF1IqmR3gFqYEpInHcj
vrklPn1kk6/kNrG7NhTKdCeq+3MZyrESYbVK7h1TlxebN2+jLFXlNibDAuHGj4nMpS3ymJAB/Kmn
BlbVHYyyrchDphMgAmyshi1vjUWBL1YeIl9urMFs5NWvVBZF3gsYHCxM/ml0y29Jr+KtHmPhMpeR
3j9uYLrg+plScAnpKjMBQrQY8u35A/89wBBwvGWCWGOQvDDI4UzP6FNiCXU7E8kwjFCYihLE/lpl
MY2cA/pnJoBr3agxhGQCteFdwpLJuX5WO+PlQQiVoCY8bnJNEex1Us9SLm+KtU5UCdjVDt6rELK/
0rFjZT4rTMnDrXkGZx1Lk8grotqc+FX0+ER5jnJujs2qd8ikwkNB5Fps8svLa9oqQMsLLPLDOVvT
5KP4iKrVaskTC4GT4ZHojrycFEhOkLB2MOxMvxAAVM7iF1VxpphWmtZ2oTvupti9tDHJQYGbeVEY
kJhDaTe6Pu2Pd40Bjsm9QA0c579g34hZmy8GyC8rG5PAbkP9Qe9csHr8rkQhIqpuHKKZZqFGbe0p
wJIj7xpv0X3QpN8HXqC3vGGncbRtIjrPeE4VzntalqNXsusiDb0ghR/HCHfvj0TZ1BGE7V2SmBdq
6nW8xjpDsL+bdz+xl8UJKE5MDbgmowKV7sLiu6fmbX6jIsJKsmLUCaW3O2xiA64v4Xb376FLtnuI
9JmNKtrlwoYBcqiPUeUtlkBBpziFvqf4hXRimIPVqEpntAdxA4K+gYZTUqGfdyXamcdTbez5qmiP
q65UVpYlY1NUWSYx4Fu5SpaWTkwC4w/hdR2BfIA6vp6SR/QkunKh7DRMw+8itXwfH6ZlU5iKNvM8
+W4KYGvsMrQxafH8xv7odQd5aUBETtRMOh6w+3r7fLAXinsvBLOlHZzdGadJ25gwqXLjLg2Jw8dt
zaNjkGKP/zKayUTwAXAzbUBxXl3iBnR87TXTHsaU8WuaJ3UB73w+pcu6qWyxsjC9huiqI9wuHosn
KEZTw1/tveTrBAWByMbWI922UFmunEGrHTrYVIi9dW98cMr7G8nUfQSR8MTF8WKnp90GFRKvrTAt
X3iFEygaJ0xMeJK3rcAD6MHk8Vf8ZDHV+kHeosi7954iMs9gtTd+vAQrbS6qRhbxg5sdb1Bscp9g
BYeu8DnSS99wQ38hh2db1TZ1ta60ZAqObcJGxJ+ltw3S5BqtV5i3jE4tMyXIJuU1djvu9G24knel
QEA96pDxywuTDGx/ud0mRcHgWNSKKDN7SSVZPuWmgQM3bOQ7EEQV+VWO4q41kL+lJOXkhyTg4OQF
be7JnzzkFXKkwTAMCoOQru1NWCNOWF2UiV6rMlCoI/TPVmCG6QqXiThu6GSSdGCeeSlO6NuC3qKc
Z80cx5W2+Qe36q8hc3dUunOQWANZVRAG47KAn1uO1a7uRWvSdIEsl4OzOi4TxQQu2qoVkEMZ86mD
GEBNzo9LuIZ2uSB1WZXJtqKgTMbps+jamKRqsnXql1Vc2J9XHFYpsLEB28HBGGFu88ooqhbK0k0G
Nzctw8JGJY5BRLRV6MZ/lDBuaPQAfnqWisNWVFWxJ/TDPNWrxAyfMsVJuySYjI4Jje0uypobTm+i
xJdlFOcihqO9oqRiz7TyA2+z0rQ9BZSp59tzwact/cO87z3NNKdaP0MrpNuj8KltOqeZ8vZJGVZj
rFUV5TRPKUZOGxmpoSGK7MzC5/o6qMgHXH4codouumicudY9ecbIL4uoxkIqlqpl9bb8Gcd6wSQ3
/LCiwMvg5P2+E2C6k6ir8EDBWkdL8+3nfGmcm8ll/W44XNq8/mbne3IODcyBklTsC5vi/9y/jn6f
5ovspjit0R+3V6QJ08GKNX4vM5GQ7BPGpdXNRNNApGjcN0UoTCgWeEDpCBQP4VA+n/hVcVWd2wax
NPHbXeOtsaL5kC7mruoQesdL2pIz7HXEtNMo2rN2o+PORqczPDWYNltcTTc6iymtZlRG/sghEfp/
WuemG3iiEk3QpbPrRIBJcushDJqQn1YfT4zMuDG1AGKXGGXrP6Hkhlyp21CzLso98rZifzpC4gB7
KBFKBWNsAXal3rd8ueDNcLk2At8NThFYWVgpg6bV0Pd/TBvWKlPRHp/DCRS7JZbh/QmPIGGeG2Si
nGc3/FibdejFjRLxFngjOelsPNhmA0N8lDlUYqLFkGczB7QrqNqil70G7mBQgqV62PGWF7n9vX84
slfhc/pLkIgIo9PGGB7FlP/zC+A1IVA+BC+VzENpt49cIfpCgxydd9u2+ODOu68SaV8V6jqBsjAv
JSXlBCvWx2aZcEF5/FTe8avyEsj8zB8y83/65JJleVPzxOWnspPNF+mPBWqu+47irM6MV0/Wc5Xl
SOMco6HM/eYdGmHwFDD5z/qq6rl+Awmqu2Nx1bjOxlQ6tG4OwTHhrzF4Maj4dXzcd/bFVWmRB2Ah
xMS0iz+ySuf0cM9WU163ZKo6s+/y2ej5jBC6ddhPp2Ce9uuni7sR9Z+A3ThxF85KtqpkKahTgqaX
sbUSKv3uWrHn24t7acDaOO2mLTyrNuYyftHNEk3u5MXp43VgQrp4845SZ02+zy/pbTiZKKU+qUhH
ch7KyUIWXZz3u3KDSkpDSPEBNeiZ71kEFiqINDBt8baSdXRYOfuC7gM580VGkmTxiHEFIgtJuDd3
MjC+RyY27iSB47QTN95P0c2+NP5VwrcUtGPxiHgRbFVKo6Z53OuWLyD1ZA2T2f+mzI4bvGOVi68H
MlB6mjvXqq0QUredYg/ZgfHGpjrN0t/+0FESttV73SOMNansEv9+TUqLEgOyCfZmYZy2P3CO//fG
V5dFPiWP1ur5gQtId8a2LdrvC79SPwBdkljB/AgYCEnbHRQKhiPDazEg95KANvB8nT+VIrAoWI0v
cfGpQnCobYJb3XRO+G6pYb04+awBUqfQFCKUnkzLvsifwrpys3dljlq9RF6STWYgBndqbDgClPEy
GcMgo5IdY45ff2k+8INlR36JwNgmdOUjdfCjD16Xh+Cdeia54MvmlWcsxPmrK26v9lbwlzq3kwjS
gOyQQhHt/um+9g/BnCprcSdrbwHKky59EUAA9abMGTDElUbKMc6ez+r78nFmE3o1chSGaGeWuJCS
sHHELNNXkBw6dYcKVgG77PhXAdKiH6XCvHCR0UridcLarwJDWWTHczxkkAacRnQFN4A18dpMYb6A
U8Nbz7zqoXJcwR6gdW6V2si6p5Fp+uVeChcj4x6XmL0NxAR5o9QY//huKXZRi/yZZ5+NKCRHwbzo
afaEOo+D9p83AaqWr2m/kaa+X0IKLxPKSdyeN4/vtu17/JkUyzY3iayKx0eKjprE6ePaykxzn0XR
r9JIq1BOkwDxREXmEtbAVsRib8niAh5WE96dHedN+vruoeJT3vXskxCuId66t73kQLk687hngJvP
8YYy/bh+irWSYP0dWCwJepiGCV29GnKv2QiaxLZ/tMhWWoOnnI/A9YO3nNyne/t+cgM1ksh2AZ/0
Tk7sihMEh/O1BDpP4K+FwAEeenJYQqWLqZR1vkgGFGyYrgAmRnDuaw1ZzWXc0zOKjomhatZC1DDS
hWHEbbgK6p8AMra7XatxwMmvuwtvYPulrEJ5csjsZTu2alqmdKeqfvgGDccvlmd8NAcxp8w4VaXC
8ETdEPsg+qwvujyzvVPj3RPEm9iI06WNXJiTdJyWyRQFfs4LEweTrA1inZ4xEifqmpZJwm2NLwb0
rBPnMdYtx/v9fEpjJ3KC5bor0U1EhH/wEsg00LxB2KrU1gse/izu6CIzBwJC7qEnMBgkSE0xTrfW
5IWF6MysgcCMtnP+/48ZiVLyXC5G+d2ub50G1zXABWiLkFylO5+sMiWoGhZ4bTyeslBBtqq4xDCj
SrIhcvkXYqMg60350AWgFHADZuBEZvgMvWEPEfrnOlKftBo5evEBO1CwENSPV/H/DHwTSkQLHV70
0OghjyD1MTL1ciLbz5U2Sf5UXxrwEXijb7uMUfjLwdYtJCBO6MgY4Ew9wgt2menbTka2uurKOUvh
WFVTzFl5lJcegBIowuGWa1yq285kT+vm1KMxyEMF+gG3Ii0Gyvi7MX3mRvAGMhnheFIr5e6P3nGU
L2Ffg6yyWeevsvnhlQfMBRXlvG8uzZMQFUR81K6ILlIG/THqCCXQXht5WOf4eTBf2YHly9gTl7R4
RIAacOp9sp+GRAo3fKOpgw2cB5PxSjlHxEQ336zgBmAFOklqHvPwIcBjEn754Am/7Bk/1ZeEetqG
pH918TrHCNU2uLY/dBKv/H5xApADrn01btF1DqIr/zJ9Z5mfBG3rQF4rKV74SfgFa+GcARwxEqXL
cKBZ+nVtqW2PUlj+BEcYfMK5ur9M5TU4Kf7kpOoUmGYifLJPZSZYRs5LliEsKffN5V8tlMNpUmSO
C+RFivlAWL9ZKc7pjo/bi/ILOvXKzyyueKylk+aXJNUc7ZwqdDRAJXEI4Te/nh5t69n6QgcNCXsr
Pj+MT5bNOQMhAiDcl7W6eayyEZRHa22AJVxBAcDlHoZP/UhEbPNXEu3RnZlY5slSfNfsj4W7HcdC
LFRroewfE+3xDlpB5VXjNGSGuZXgHz//KD32xa3IIOz/4Y+qUxM8esPDqX3T1QOOOU7rDh4GdoRy
rWVq/1BrS+3+pmMEksoz1P8m7cbcQsaiYxx9CMom4YXveSmeUYTTm5THUet2Ls4GP2o/H3+Gsh5f
KNmAuDiLomiUEjr2gDqOsjbBQI8przuQ4U0ksZhKnGYcUmrHi4rt6HCNcKEIsJ9zU0zZrIoY11Pv
1uJv1pJT0qNvzolttaGBqz99ESzmWjVBOPAZkGhjnILVdui2DQLyupPfuU1oxw67k8v4ikkgiBPS
xrjtzb0uvYb1aPkVzfQaFTojNoIJ4EM9hs2Qu/h1DL4RZz5qITQOFeQNOgvvXYO1M4atSKjaUbR7
ZQ47BgUGveZne6J2aJz7JxbuAjGO2goWvat+7ITP+d6WeUaw8nZ0Cnn7K1e09OW5MMLlLFrphA1B
bPnQit12ty8G+uuv3sspISqVjWxHJCopJZUfw/dhNwX9AjLFMPoGhiKB6jniHd4OHwU5nK4spZmK
V3B1WzkrFH/24Dj2UAKPyAbzHY99U4l6NJKBsA2xGHDc9QuP9j3ELRf5JEfXjyHt/S+IaX+la642
AFYpLeuukkzabYU7b4Ho1DkVKGonxM06I79ZyzxvI9eoJMPdY3wA0fvuxPpfeq2ecE3ApO3l25GT
o86CwmWvbVX3nm6pELj6781W6C8TM48K6BzOgvHzrs87CbskyZDPZBSNUUJ1zJobRVMk/BZUHbeY
6bOCjvpG2loDsdBxbgPhg2NCS3WQTp0qkokf5xcInlyWfbmI06A7lwGoaGI8YviJgwuPxV/idWwu
MYAK59bZBcX19iQ0wlM8ADqheGBSW8peHt4fRqwiKCmUq6qXxmk0CglpI8eIqxLLd6rh1PAYtrek
FxMPh1ihMVV8+9nDf1Z54ICmeTn9pMFNd8LTJZ6Wx1e0gBw3KBCWoSN5bmtMAqjicFJLil51cAq1
cCfIQ5Q5ojLX9qev5z+S1hxXTI/13q9qUjtXcCpGCqQJmhXf/07efgusbRCWgOf6Shn3Y6eBMx2k
iVZmYem48DuimWm1SFYOdidZJ8BthWqKP94W+bNc/pyamc78MELkkqEN/ALASLn78mcw3yE9n0Ut
7pD1N73gJgjqiGnVXhVrumrNBulWVVtRp/C1teKjJZ7xxgpaYN0CQg3cCL6Gl2PGYvg9H5q52zE8
AaWHFtyLJrD5Eo3gjS2bR/0/q8YeP7d540koej0zEbDDEU8GXiACtfyqAGFpcPRivkIwdUmIiOQg
6PjIHyXkCQFi9BnyNwPrjNIpHI8AuYhQAuE3NkCCInAUbhhZdoiclFlffUkzzCNIkqQ7QYbdpJXm
/sGE86rPcQBusf3D3ucefjnIy6VIcK1vCfAfMt9TImezlXlY3yxFvguPDrW1GfyouW/cUZBxskBr
O5E/nPTFzcFtq4SH9ebwXD9OXGaFO75Lb6zK2IRczx9i+frYuRk0AP5dus8XuD1DmSx0qCfLmjeI
qXDe13u7zuCPMgEXlC8IOGynjZOznrf+cGVPKEZEzbtA7xfaSTEg9ABtcM/Y5qUXCx6j2BKw++oV
FRAA+Shg3EshyN5B4ntNzCj2gIDILOEtlnoWG9LJ+xJSLpICco+hE/EZrOwF9rSYKv3hF8dAkFl0
5kXP2JiuBbLTcL9fRkp78T7hl4uZmdvws2mALB96uML9CGxPpoKqPU3/t1xwVKa1MFhKcZUQf0q1
DFozHVCey3ZLTcfuKColEYDGWw50wmcTRM47XPr5SuYaCpxC2eQfmc+fKHXD6y/w6sHMJ72Mk4C7
FbiRoFDHuZLjgBIUjkEp+MIiiNLIWkaPnsXaAE0Y7izeUkTI2gP7ya/Dtg3gIFYBFRMrNBQFcEmk
wayIHcpu3zmiMSDeZ2iG0D7N0I6MM/UCFc7JATxziVJuI8Pde/OaRrQtdQI5ZkyBIHpCDwDvGsQj
Ij5K3Ucgh6dtMfL5kK/6RVq0bs2Ao5lyRYX9Rb3O6YeW+mdvOtE9Bvwdw6BXUQ7BkRc9NB7RJ9l+
Uq9ejPJxh20EA+RsJ1ciRJ9D+Hji8g3qZ3wD3swAcEWi1Fl1cHngQLvet1ZNRGPSrwmmlBj1+nT2
Wyaazo8hha7ANCO7OgcZQVlWP2cltig8Lg6S+u9Bdq6m8E8+lknK4QHg8ManbDTl95x7o962ix/8
IbwWtxneqSJ2w5HahkNIQow4A8+tropkVVaAi9mBEITRRNP3fcrW2a/pNWyUY/KPRX3hLsNA4qtW
KyvLR4eMD0YCMU7otca1dAAR/nKH1MzI+l0XyejpaOfudcN+qt8X5WO7C/aYz8zn+hTnkH6uROSZ
5KOMra6Y8Ufzrsi3zJmhBn94qOOYgM1q5hS5cP/+20yTrnxrickNXXKEbfGnJP7km9lLwBrvyUaK
qIA28rUkzL60e/Eb9RWuzL/U7AVk/9ySW0PJz2DzLcNmqHy5yhLtbN0hJdCzcG2lnvYqJIzXBml5
jbm+Ripu+dsaSMOAXt0ELWOL7bgrMXQy+3KXB822vSMULYqI8YiFrf6L65yX47PLjyE1oR9lm8wr
c9SXKFnJ8y34D8lY/QUNSl6+iklRHlb5ZiDmtCUtPgN0teoppTLc+ZdeLjrucHoqcdP8n87lICCd
fKeS2ktTwpS74SArTEvjqIcpCQF/7utkoGB/6VlUqOzBhMFa7Y/S4UQDhecJ51qFAfo3QU2VbTk6
rt/XQO4OtAA6tm3pbyjtmgNzYnFO0mG2vYw0Aw8iwF+Swf7udvxP3XlfM4ejGkDtAKdLvJtKB3KX
A9EpMlzNnktocY3u2OpQHO3Glh2mhpswf2wKXKVSg79baVOhAr7vWwcoxunX7DLd3F6zocvs27Ie
k92OagDsj7w5vxEHbfLbmhuGDJ6UXfPh1c5oinwVUVvnwtqCrUeNFSeLaUM8ZWcGntjDAHjf1lir
NnNORLuCaDXfcvLCK6wpU3GeZJm5TAC63nbFXmot4WNROO5QQgvaVZ5W/FuhcFKVOcf+dEuX6deC
fKCpdWylQBzsOZBhj7cVXk8KBk5y28GxeuVPzsnpH5a3I5hbE6eS5oWjw1tYnB7+zM130dis0t8o
/wRMaXAsolCsViTjMdDJBJ1dXq0Ghba2JpW+mdrjAX7bQ/h623VAa9RZkfm+gXipZzWyAYHsqHXw
y6t7e0e69zdLNsFPZrHZSa3bHJK/+tJZvSq+ObbTHc5D3P8SLNa+jnnABz189MMy0mwgcFSuLEYu
nD2eAK/He+sj3pL+C9J3ikCZoT3sccujhzSNpgkL9LzjTBjNDf9IEsz3GAsu1P6G2bDp0YFXWZ41
Z6JTkFvssZLqu31c7Nhp63/Hnikrsik3npdxi9Xm6W4WGdk0A/4ffLNmNXTDMlKxMTZXvYZuuVyp
6ors0JrOcRufZekf3Q4NQVzAWoJaHQJ80eOMh1LIRwV7o/QYd4M64pOfv/iLeqDSLbPyN0dPlXi1
EZXaeG0PQORUTMOuPEdyOxkTm1X3DIHmJe7VpnRA/krJwZe879MUxd94FLSUdJG1McUsqTmdyqij
NjroNcJAUS1+qwPAUL6Kizdf5NoUQ6YuoE263bglDLuKFBgQHeal794emfuKv/udYX85f5kwm4yx
F0u8Tcn4yEWwca0VDyGocupTSYrTjaFshAGhax/kqIQVxqup6p+Ws7DWi4fX3ma4cpggi3BplN0C
F/9RRCiviOmwhH7Hz3nn1VgB5jDGSoEnYb8yrwWvii/tskz1fNhp5V9W+dSVSE7p8Dj30JPicAh2
x0Z78TI7HsAYSvlYC7eEYLbWvssPKog3sHmyZPjm34QuzdkBui7cAhc995VZGtw0NpyeopknuZuo
ZiyicA7xeSkTBTACAvhqP66/f7i/RV3k/ziU8JRXzesAfnxjrMgbguA1zlC+AZZEKkeEcW0Q8hja
X2O4oAFqGSZSyEy6AkzsSsXcpeBBPaJlWkGXdxeLt02vIFcwS7aiJcICUyxrZ/mMAjJ951eL7b8R
LnJX5Og0pKjOdjXQ3fXPshnTHUpvYIpHCLN2YRYqqwAb7YsRHV7AYirf6PpRT3Oo8/Nn7xHo1PTy
1UdxNm+R3yBdbeeQF5C+5laretuPk2GNG06V8SXmvtdBwyFitHoKMKKUsafPUDhSWcxWylBlaqOP
LuJCa4nP+h3D085/hVj7HIkMTAn/RUPie9UbqdCKcy9ALiQE5wP4ihyPAIKpb0US3JRx3SGovsPK
SOzKkBgOjCaU/tjlv+TXf7M23ZTaIDigOG2oOMNtV3wA8alwHddyWnYeiha5tT26PLIXcCxCLgZQ
z1qQErpcr338VBblbV8qjk03Rp26X79HgR10buJu6TBNE79KXlXiFGHshBrbXFzvQRqlbjIvpUBy
8m7L/ygNOMoKJMqvkhLOPk4Fl3U1f4VSZOofv6CP1zJTY6mRgLUlcOive/t5W8jaFsUROdz7vnUX
uOh35IB2kM6BMGO1IJZ7DTa7K+qQFlm1E83/829USR3kJdgDj0eWJrwB8NAtBQzmAK2UQTROxI3W
RT95c+v+5RXNAseL+Q5yeWHVYOQ7Jub4RR6qWPrr056Hd9AHf2vLMGKSPzozzxWunGr2XNHUvNC8
wJdxK4jx8n5RdQzaGTfE4lUDmzr5ZXhzHylGAvv0nol4309I0ZYfMkJU5jPqlWA7q27DTKOCkBIs
GMadwWMx1DthmmjmMoUwZ7cKUJL7GzDfb1MWbQK9FpuilimghO6IpyAu99m+9bhzlbaGEkiuETEd
S9kHvGHcPQL6Mbtmc8EeId+fj0cd/fU+1FJb8S6o61XyCyJR4x/B0Y8NcThqJz3Scbhk1hyqeNmq
A72ZLGZMebkHQ4Os1eqUFvD8nFGmjtle3wjeNSz3umG/Z1kM0jheHALFW/gPe/XZo9rr/e9zeprq
0BzAyxy8r3C2fvlhTc0HVH32ZIiWuEjV/IuFao1DoTRHCfJpt/lv/mphBLaKGBIcO/eVS5A9DpWj
wuE778FvZZkcSYdoD4ymGxMFPMR9xs9OAp8dBxrH7FEkksN5oKIsEqC9b0kMRw6uWc02oknycckH
x6wgHaGlpha216VZYIdA+W+QC4z0Gt0vWJcd6Y8Tee6I/MCJHtcsP0Cch7mflVxxUY/kSBGe1rf9
1QafduV9HrgWES/FBzKp08X+pm51MX9sXcWNlbC2y444IDKFx2zhB+oT/Wo6L9cnGmyaZapzfweW
b+Uz3b7kMeUsrnD10qX8HfWrrypapcTurdYjTerLa/3VMyQ3KqR6ivw5Lifykok6U1AKQpcqRaK9
GK7/8JzyrpVzxQPwWLDOMvP9PVuBfudz+p2yTMq8cNawhxcdwh24T0pa6hwfJDQK7SXzFsT0/WyV
A/+XyxwgsRL3H0+jJP/WfWN/ziQPxoLQ6ryd9ao00CAhMib73ElKuB/CnAPDML5FlXuytyKRm3fT
GH5m7FkW8SEI4R+b88L9utcFKg4C/FZNxcve3GddYMmo2OVGh9k4On54WkooX8UFDc+Nk2X3ftRp
9WPh5jSeghHmwkLTCq+h2N4Q3yxkmVoGDGR/HM9A5E25u2M21gQUHSy1MGHK2fPRgXBFWnWY0+Va
E85y2quNYgiMIPXrPyA/blJEwlAp70HEw5n3uhJ+UMdz44ZYdbXZTs/Y16GrHArwpVdPYxRqNGPH
r47/xgqWaXAQbmHUZDSg/6lpalnuLQb2s2Gfts+aKElKtSllg1hXT8JxvU4nzuGbss+W9z2D1V+2
gtH3htsA0NGWWr/RuqjAFUt/S/3D3n+zQD2BkDtCkYPsrvaDXIORPmw/yKhX//yeZ2ojzg+QCJJn
29PrfAyCsiQp0aFkkMwXQ98RBVnJIdgsjYgK/jMDb5PJZyRMl6WEuMtis8/FYkWGMHUSgaRqxq1Z
EyxIe1fFcOXUrAbwdrTAXVQwkoWipdZCjOokB3nj8fery9RVCbBMx/+adQo15g8g8QQnnq+xdASH
8dIAVp2nGdBttQ+GjLsTayzqH3I59xf9RrqPZFTyMUd0VJL7Ra/nWtPvbQ+moy0zbFZ3RuYUQ4KK
w5bfZSia6pqOXy7hZqMmgRQxfoU4czSikNYEeqe0LUTWd0ODuOaFrSVNj4ynp37GabmPRCYwaekT
OPA70hpT3utkpKc0On8gc7pciW+d0/aYOw3htBzE9tje0MwnodvIG4Sn44mH+/96t1JhcbWahhEg
M5WkSvrpEL1xxgtW/IzGBAr7zw4tMG+wGL/JDfZabp51v7KKiMY/hY6cOqGUaG6iM2CtrTDCpZIn
urE+h/0A1pTkLE0RyHIP3g9ePSiaIIAuRTlRafA+mDTiFsX+q14RyyCAhq9mkQOKHpGrQULgXTsi
bti7BPsTxh9ULT0pVFv4iXO3A48VYVXjI3wBc3TqJCKa0SeW0JaB19o5qAiyrWdQqw9YD2X/+ywa
ku70koTEy4+qA26DsUNXbaq6df0+gZES6RT2p0hEBI+OjOBrJNUE2eIbOZ0AZSnlWdtLsi4NwiY4
uknICG6KOhmbWVPmrIsWrKEaQNTbjEAz2+AVg1M+Ud1c8VCGap97axpol5Q7JKXKip1fvcH4Uwx/
hLRtlXmdVDhu+K5JyonwgCzwUZMG7ghvhmTZeHtoqmmh3sui7VF08F8KMQyD3mv2aME8Jsw2Qll8
yjJlCtKSBKxIoQX/3zh90k3k4+5IcNKtpM5vlRwl51k2b0DCHOP3nlWecvDUvGiLo9+dRq6zs9gc
U7yxdkBjQ8bLKZbY76mTFvGXvJjqHXeuZl2eQNN044ctz3CjyLeBHAwBPx2SxqXiIq7VYFe7SH4v
sRULDEGkhvVlM/XggMG9UfQTc4ZVeWb0q6JFJ1zS9DiSfeziORArTMCeYRypR3/UOal7zBCN86RC
gMA7Gb/eembsqQsw1jCKwHyqJTfSG0747bisHOzcQ38E+4QmQRNaa9tEMbEj3rUjY9r97QihFM4c
cH7U6KZ5NMqHT5MN2a6jrBRSC8RQVt5vHU9YPZESwKMdgGOBcsnVFdRcpXon74H02Wre2jE1W3tB
yyVb9oNIbCG3iQKByiwiazFCgFwMtWpwnw+LDmUESygkXSNovZiRJuCev/MB5VbL9jmljhscDnIr
uyMONbHcosQJGQQ/Fswecb5Vu8mASOMx2NJptipUvEl4p49Ql3B6eJCsc0x+2YuttzdI7srYuqQH
fTJcubxOxvCHGKt+k2tQuLy+kiIM5ypvDQuuhQoLXy3oLxHjIbMGkgrrBzDppbititSySjneIwKI
0DxkVG0bLgqY16tsBIDGHwLf4zse39hFNk/Krx1kvk6f2H6c7+qtA3C0dT2iXGsjcPAk1TjTd9hO
m2IhhHdzV18GNVJqnAd7ahcRmnDwHh7PWDU06BoJZQt1I9dzG+RuZszlK/TVvt5HQw468jQKCWII
4Mk4/d3D6W1qUchgmbkn+nMeDlX7rK3vJZIbX9WUAbX/zoxsd8XLgqmGaFhKgbthOYXigIoO+J8B
S6GZTAV2SA1FWNTjOJnLR+DwXd0QUPBn4CqauszqHKyoSpuvJ4o1KMqcn+hDAzn71JE/MDUcsIm5
Hy/ouVQQPzxfSDtN8P0hLX9PZ0yCU5L7Mr5ZQDQR0t6vV+auDaogtpgPkVXUSrgXcBjZ491wNG3C
x82PE9zbsSAq2JavSk3sAPAXzPjqkvAvLemDcAxdAJXmxl75BlxPGVO6P/Ri5bXCLh/brwBbGB2l
4hQCBHI/4WvJbh8DkDGE/7+yn761g59bG68Dm8Hamzd6AfRYsoCeHfP0u0vpRQ4C4aSowlhnTqBL
nQkzJWb0bvEwO62leaOZ+LGqhCP8WTibbl8lD6N4zR4IKqx7d0pUi1qpljk2oSRxPKozQ89IdQU+
xAeKJ4F4wayC1fq9Jwg+Trq0hl6gn4SgY+mPth8Uuse3CDzY72Nx7Y64IkTHqbK6yCBlbc5VXgQ+
0Mx/sGf6D1wTTtxmgiaYU/A1/y5Atu6tk3IdD+d1EUj2Oi/q9/27KptvAKCUjPlXgGzyn1LCybKM
EsEorhtnNDVlAJMMVgRv8EVQrcFhv83Kk1/xTpIgOb3UVd330MGViAAlLVdbtL4ON3GXXkffTCRt
0OjPMytcQKu62Ur1NSO0zYtBWd1rR0IsDyLZpvtvgekomIgO+9l8vm25nG7NVLdx2CoPLO+G9Q6y
+qUHepnWgRR603epxIpRXtgnjxXvG3yCX/uW1EBa18VGF9S+/rr85zqUyLUSMCVrx1mSnxSmaU7v
92Mfige0k5gEGOptzRk1RnCFVgXpOAm0mx299AJYszlWICKDK88jMvqa8LE3rZLzE+QpqUTX+skO
2cjfbYNGMpTnmYF/LXkC9TzUSIoZJftK0aFN7MqWezCZYxBEpQkJ7Rh8DfUbTORoy/wnaoXJVzAm
yp1Tpq+rt7EX/tctNG593Wt6kf4As83j7bgfn8bx8TNVDiC2Fj8URBVpQfnwx8/Pb+T7L4Q4dij3
V+PCvaPADenXMFC32nVu0iI4ne7Nd6CNNri2z+YVViC1+evECm/484io6Pa8LpLkWHjAaxJ6Zc5s
PaZvXJKY81t4eHsK7RVjL08rVQmojibVGKLYojTka+5Et34IfND7ZeN4a1+fopQ5dZHboUk+MDlx
N5upkP3QBeDl/tsQ/CQe6ieaLe4kcWsf+FOZx1aOAHkRqFOyb4YefZabf3S2pAiWhhOrespcYEOg
TsNb0+GUsz3cfovf78aSUE1Us6ymC3AUIRGnYEtFA3k7D1J3ulLTyuQuGhQccebYZYuq/CTfvL2J
jUvB4w1+3FvTiILrI/QkjiVLAi5crrp9KkLI1ZA/T6D6xTH+mB02cnWXlybLzsTygOkE9TWLEh5S
3irVjtyfkTyI5Nj/ulUZ0CN7fqHX9pyNGBTRR6355KCvFYssf5X/5nF3Bo1lUe+kRZXqrSJJt0KJ
Gmiy6hlDsTyAsBXtUHbkExjE+PocoNAoJjMptdAfE/Ri5WexhTWfnzYr2W9XqlXtH5x3Gm/6dWte
mcA7owMsZavKBUlXsQLiTUPI0B/7is4UcgM3Qm1NPWxUZadDfjy0HjxuLAf4eSfeJN3igWOSXxI+
S32drxaWGCKEtlNantsGUGyHT9lSGqPxQuQC4mVGrAzSvpj8rzAJISrh0LPN8wRozMEmVTx4NVTv
zPTa3FGBGdlGf1VVvwE3KBGZfJqG4qwxHggDiuRYCmVubsgaQ9QdwTpt2b73jf+cSvJTT93sYrNc
ThPZsi13n1cEiJus74Fd4POjtpf0gb4f+Fr6W+uQcWwI9so0GU1u53h6PEktmI7IhLM6HkdkZDGT
wDsbfBrthor8y5WIayZqwbCYCZuORYj+zakXPMT+qe5vg2nphDunAs4UQuQiVUsH67f8t+mPmiZY
U9E8bYMH9sdIk2W9XtOHMNw4yAksbg5883oyq8odinwXGyVsAno9C/i8MkxfD8RoNHxqloKhsAAf
uIbrDlg6qrAcTnf0F1uGu0nIrMVcXgkAsR18fVMwUaYRYOv7WqlorN8TJXQtJWkHLd24kKrcUN61
7rkNYEgOn3yx8CN1ejk3MrhqjrDoNMNpq88e5QUUr4k9OjNIXcdup4yw7KqQN7jyWyEmey/c6FZT
38X4Iia/1c24Z74Jfuq3cze9XTpTRitf6ovDvGqm2S8pCMHMC6UD53mxgGV5xxSTyR19AcZ8PJa0
YC4/luLfnapMS/ukdlTy4Vg+Vo34Kqsp/Y4UtGAZua1gRlf+ma930+qJ8T4j0MMVXkKNsI9D7bw4
WaUCAcWdeOtF1ats0WIVVf/7l+s9UQK1BjpvLtVSClQ6ECume2aZ27iL0PkQVMwGMRNNM45t5viK
aXJ/EXMMW6ChdhP0KXt2hyoHI2ATS+Vao6QNC9ztmutJW4O9H81c7Jc/Q9MnLEou9h3mrjvn3rVX
9VXs4kKSsWkLZZ0bpp9W6IInY5Kj5p/xtjrJGZEePKjinZOvldVHHHjDrjUlCrsgtalUD8qR4lm3
xZNPvOSOFyufeZJLUYw7B5T5AOzZ3OWVpsmGO69zNWE2nZ8QzGvbn8D3b/E6DlXqBr88/ikkYDel
Y8BS9rpa+25pnrjNSqFKqAnoDlrre2Hew3C41k7bpatqSfkZank1Dmw4OKMNsmsCMlS0v288Uirr
M4uOmkS/S7wc+10XBPdZs9MQK49Eq1WwtoA9JUBmXyejx0Hibwrk5dSGXqHuFCO/lCrV106rRaHW
a+eJxe7UiZQLS+gI1uCLeAaVFLfKZrCyJv0SO/cs+AQAv9SkxQHPn8El1PxQNGPp4B67dAARqhep
l/RD/DDxjMFIikRZEJ0IIIk7LFywvrUzQyor0JTs8KECL+/ArU3vW3wNzkVbx6NFDUT89Utjzz2d
ZueTqQ1ok4b6GM6il7a5hvz+w4oNy62sgCYcMZ8D1kM8KCHnzWp/O0jcGmIwpftG6o0UKtXJo09z
AESf10j15aVBNHuN40Mj/nvp/wnLf/rQ4SynNcH+yvBWkebdiZDPHvFaaEMgc4TqylU99GPLFjSC
SEBHRZedJPSIacBXzbCK+OtrzWLMf0Ma66Coa+d1V2aVAs8mVnsqiFyC3J43UyyWxpFaTBCa08jp
EJ+ytpe7QvHm6Fu3OjLHh1sc8H8419A7gCgOlBG12oBQYGSCZedmPqmhLpMceuunXKFyoHXb46Qi
+0W5FGV68IBYwMd8i73otzHOuknCI2Sq1qHoiWcXG1R/XSF7y1yQsLP7sJet8b6GEj73Yu1T3QXW
KOsYTA2iclJ8KUqJchYJKYpgRrsXhj3RUAX035cQ6owe8cY2QuCPFTiDgHn3m4A7rQluvYi8J/mU
5c73pQC09ZGk57wd4sR9DIjEx2OQW1qsTcEfwHEdXoD/nZsyfAC4cOEicgyJn1FzNK8TV7YJKiz+
vOmDhZLJBQ95nITxe4gCj+Fxy8G8PUHxXBcAo27Ld3xP0YHfjA8eWAjRvo+z2oXzYNKTxK5V1HMo
G7RK9gfcYvTRwj+/rrSW9tTeNiJkf6+BNjLorx1mJG/8wmrHxw+pfn+6nlxPtzZ1ov8Fd7ZuAf2p
DIfI4K7wW0QEHoFgf7+zCCU1JmMe5Ytsx8zXTpombBihZHnTvEyMsf0aLxIltWHVsRM9ir4F2Od+
b5uk73yW2fTB7O1SVga53Kk0p8hGrxlN02RObFaoAj8/jozqWYn8LiXwj3llQVJs9mIhnKHxSrns
a1TIfktO2oSEPZv2wny63JmmMD9qCE2LZUgtC2ad/SFSsxeUErnRMskfCk2RGcuDoH0yCEVPtkup
NwAEfJCilDwfXcvxuyPfjMITGMrpLDKQZeqF1r6wXz8dRdBABt38kUs+V7a0eFu5xFYrwT6GNczn
pz5s3+XdJ6vWnNIZWoXJVAj/7YxoPkYm4d5YEA26zQlUzbA0x/O/wr3q1mJ3BkXjuy5ENr3A4XOJ
sb4fUyl/VYJKI9Fm8uM38ajKGHhWG7J+VR6ySXNNJI7pm36cTJ8zk0oDMN9SvtG44Kxc5NGbdKND
Kuo5FbKhYyGp3RozwK2w1R9L9/xmnnjDZyoIfjUl6PIPTjVi5ZYyWYRenKh6EWhUgEdboNmvdaPQ
RosH48Qj6UY7IhR5d7PLdevNRGy+uy9qtoxSw5a3Ga6nCNGbVdUp8W+PAY0iyqjLfKOpfethI3U7
UUPgqASyYEuI/bfE6rpAIyPmR6lB00ZSsQQ/krmaFVEZoYFCvZZEyHV9+AB+HdwR6fZCKGJX5tJs
GhltXsYMtCzl0eXUXKdfKrHf+uUjbBJ5SqZj8GBfEhZUG2u2BdiV4ZKIVi0XVmdeHyFXoug/mAme
ydqBJtDRoiwaEjD+cIL20XC72l4vTc5mlm4p3IUVi7gbBtQWe6g/+VVMO0e7Lex6pjapybfjeBnj
QvJZuJx1NdqW8+goNb/D9gQiZURkPaRCkoj05gF3kpkNSlzH/MkS/4Ck/1QKRQeYT6h9LkduR1Oa
QQstcqyIvQ9do5jdr6/fsltMDuewFU9YzJ83VGPRPGyDlc41cKwa8LSy+yss8EjOX6EIKQgxoEvd
V932RmlabMImhT5TrNLLs+5AVuCgqANoHr+aCW8iaMTsykUHnGYbQlAGNIoe4FZAc7PH7DwrXi0d
Cu/QaVijt0rY8IwXoZwGgudsfNXeSVXuTfy4iuTM9y7s0ZdUB1DT6ax/cVy8Fjg1gBIk7/XTH/21
1szoGVS95nU8zCc/2STDdVTqknuLnFqM8kD5+a/mLzAYTkKkfc8CgPnPR5QlTBPIBfyI9OmwgkL5
lwdfoyJQzMLgFW6RDs0o9hKiECYwg6qrVKfCWUamjYAuaswAFYibrP+YQ7UvF8sIoynzhsNn5SIS
URL8erSV81sjb9YCM//zjksvVpzcikozMoNq11fi4i4p7eHx0700IxuoDDMLG0NWAhMQ9kZ6QtMi
UdF17kjjDtxFp22fcyiEpI039KFsf6RKKC4Nj2SzEsQ3JgXxSeUL5vXBSoZK0mx1ldxJjmTGI11E
BDIvfx8J4AqhHfLXU8G3HhUCQnoP71MwHvh1/E0mxjyuKZw3hLiVOu0ksjpRg2NQ7VhOITHtp0hT
sKN9OXxtkjzdX4YAP5Gz5DUL0YQs8CsYL06bgMFLjAlG4tgGsDLXEGHM42zRs09UBStz+7+pSJsu
Pai0lC4GjCvC3wZgBRNWQQ+UidPpDrUzr38k2x3NJGZqwgZ7lssNQ+Dlmh6YQpTPug0Uy1sEKJzU
k+TZH43cAO51j0kFAtTkU2GCsrLM6/Gx8RQ3AIqjv9/Fxkclu/cIFU0Z2cr3H+CcaD/232TtW8+X
NwBy9UkViZenOQUwDT2oJUq2D3hqwS1BTz2/XIMhvvcQsIq1xbjxX0t6mLx0nGCjDU+wAuFMhuXp
Rkhzq5Ul/XTJJWy1GJRdLFlynSjeo56mRqdmIuzsFdRFu1SI6wbyJYMjxRIgbTOhXBHLePTN9MOD
VQQY89rr76bS+zQkW9ZLnmtnN9NnZSgjJuBI729ww4Y1NQIbx+WYA1KpEe4st8975+kSYwNCzMnO
Cl098gi2Uud1f5J20robvrd7Xwys2/Nw3kGBGiYe/TzPNAHnsoHby5/vPHZWFzO2HtQjYL6w4uJI
e53n2mgga7J7zIZ3eq/fOJP6O4qugZCT2r4YF2mmQ7g6IVX4ZaoUHblBAQZGhMLXmSzF4H+tbtWP
WvX3XOcH2JEdspyRB9mErX6uxQ+6OCOQvj4ckWnGMkU3w/iTi140gTkKIGaykpKShrhxywXDPIVO
HGFl/2ihZmWgXIHjAw2G2YeIuRLtZyjhmpxoB2hZeT0anbDdBWLIq1H7CfleKaDRrQMfUFwoWeZB
Q7KGFCNHRw9KZgaduNM+XQxn1EJ20FIER6ji7uy2Qw2dbT6h9qg4owMidwcdCb94nLperkjajz91
dNoIRX4Vdi4Gield+AZ/ziqL5GY/cL8J1AYerqDqPoeGb26rOC019zyVeofcvojWgE4PP6Ou2pzH
1jVKLPRPbEUfMsa8U9Tlt6VH3W0JFXlpr5BLzV1boQHAWxL+KJFPFz7cHnAeaIkFhReYuApZILGy
Owwuw21CKjMie2FT/q6F0mDhag3JbYNva+SZD3QaNfL7dyRLT4WFYl1Av/vQ0yR5qUtSn3KCyr9J
hRYlOF8YIcyClKmXgc8jvg3OJYls5DdRqNs9D3m4pk7UF10zla9IiZDFJYPAOMfxMNm7n2WhuzN+
jI+Zo5lUwaZjzhUhIcjFvnkVcJQhxNysWzX8p0CnaJjDbYrNKKg9l1WYyTiSj7dCcPFBSBp/u3nG
LmEz1jvNJQ35UZGrLvsvFpJ+t0BPKR8fRB6B8TyLfOIM3wuH9bO57ZIoorYw4L/mg4CW8ufQnuUl
1i9INZxQ+HFv2nNdqMXpwBRpoVkHdUfJrcckS48cV2gSfMaqe/AliHp+SVvbn1bdCQvfQaplBw/m
U2S5iEhWRM8ajBV4x9Xc1h88VmUdiBEvJlLpejHXTEQYyeHQmyqMyLyVmLZsxiJmUkSWOaKyqZOC
clk0oXGDr09JUHMANObYALMelw0LRT4SXJwiegy/50Wjw2Oz4EgGPp/5d4Qy1pt/7tdBjDbzzN1c
KwYGMZA3FHGvApWWf74TSylMNr24eYL6vJaf7b6xOBjtUY6HheVm4HT2N71TeHoE66wg0X42Vq8t
YrV82K9wK5IfG4uSX/9Uv4JYEz8J/wvryyyLY/wYV5aJ2aRT5GzNzsmOoojxEyj51htpEaCzygtH
MIG6WyuSrPdK5GIW1sZNxZcDCuXu266b0wgGrvAjp43DRTA2piqaIIJTbnf5382jVMCI3SgttFXf
3eUqv4TKufgQj9IZQSK1xs/SrCKYjDFsDDEobUQh3fgRDgcrYewc5MyvV5x2YKz2kg9DFFzGwo27
BVO8/X6LY9eim/ljQ35ZKVxBofpCNeGtJWUHHzZ1sUdnxaFQXEisTD3ezlncXAMecVyTz21UL//C
2WpCgNQkdyRIyBEDW+J1qPyPxZn5K3Tvz5h7WTGCmQKPp6F5cGfCBhh8C7E4cp7lhrITpNWSK2s9
GRA1vKI/L10yVFsV3TXLB2mup77PQutJ7NCycKCXwgfHwCPGz2xUF+6JgO4vqZsV66yY8MDdeWlu
shcvunv3yxbBkyCykAS77KZg6NqybXuDb0QCfAenrnr9n2sEY3cR0r7yEgOlch8dphVIDJqdtVLy
wCdkYWjbo0PuOzUYjUUMDZCOzYbGTWY6zRbJ12dfR1rCiYFOEQJP1NSLKFa7xTkYz5F89ENhykE0
lWKK+wOyYq1StMpK68ChvF8dr3iruPLqqaylQZk49UKX4Af9cTpMBasYyAtjofdLhPrWkpc4u0Ly
F/YsyQSbMEpOraqozwEQ4lbDsTBo7iFLB8EQamb57OuqTceYU8Wj4nkyRxTjTXavPXcbBYeYV6dz
GI7NCzSyuIyrKiu70YbGd/PZN8u2zsvduGRskcHldhcRqRcsHQy0VOqPDWBoV/B11r8vz4mdW6Pt
r5boXmlv1N+cr5hx3AUZqlQ6PHd3/pUBp23ldQKvowpZV3j19IUFqrvyRxyVmhbxHIGxJ5ZstMRS
dbzPEufECyO0Bq4IXtZwGvs5Li+yV0A9eH8lRV477RiMhIPHCuglhJChDSe5ByjbmRyAMGIzYu26
ax2PdGNQzlbYKY3LeMLGABIx97YtXvtuJ51VjtT9Ja5SkXgaAFC5lGxVKqnFANZhTaY8DsAa16EJ
DYSymSgrHblbnwXJSVKZAlwgqeBdJPgUqenIrdwMMBe0+oyebmgjPys6Raf3xg5hmolRKmndj5sd
QO4hk8F2TZziUj2maRYk29rNMSb+oirfNd3mdi5HphijSQm/ka0UhAiYfpiv+dyIKkQ0t2fJCcVI
dodrtJOJgtZaidW3VKbjoDOBc/AhZafc/Ii9WtU+7rkvTMVHU3z/DBiJSlG8ffeLBqd9vYEQqHmA
Gq0Kk65C4Z6F4IgaBOLqRpBVcw6ihqBQbOzhHfhn4THqAm1xlKrG2+QESuRNAf2X+mh/1xzrNQT6
aRdBa7obHa4al7VhbMNpOzgH25FWNtcdYrVKy7mCP2+m1NmcSrtsbwfw4YAYlKQcdXv29PP7r9sb
TrlAUzKQYvPlUtMp7SztDbJozJJW0kW6mjVupxQpUjQ1VdRtuB8gFbMA0F/m779oIsvcYZVPda4R
0MO6JXuAeFcAmT3835MMsnIGmpiJ8CPRurHF4zOW8y5fYgvF2OLbts3Cconn1RsjvWUXs/p0ltxc
PsMdE4qm1Mv3wepb1ud7P9YAcA73fcmZ3IAPaUnif5gPvf9CBLSYgAEz+rtOg8zL5fFpFgpjmbXH
Oz+nqJ8ZrDTAtiqIkpVvgTvP8zCY3PYChOLGUi59k5M8PWOQwLnyst96nxN8ULhfuIR95kZHvzZT
RWHiRTbkL+03yJMr0vOk0iPNYZjTTDQbtc2dKz48AdD5Lt9os7v3QJ/NJTbw+VCY5aqpdTs0fXUO
6ORkEKJ3PbPO97QDtsi+X28LwyVeIBKhdzlt1qUcF8Y7WViQXH1huSucltQjXtVDKOVHkWNJVYho
bSR/RAIb85dU829A8KBkbYsviGvxpIIUbAXy16FvLyjQuymC0dUDzPkbw2r/e+GxBUafTCRM65pM
DEcuCReoXE7wysTUrTflsbgn3vbhHjVHNiDgB/6PeNvR7/MlnkLBDt+be1CN8FcNNnTcDV0Et6Ws
VKaYuFB27nkT8FbC5zJVOWGJ8CLY2w73jNYQSMdsvSB7/pweoXe+/Ng7xePSCOqHD7u0rnJbxwM6
STRMb1hQEsq6B/PzVvh6VJ+fPjQ6Jx+es0KaxGSXMYbf4EkzgqbVmSo8FdsMdOkYOaxUDShbrw5H
uFGozHkcgkXFmxN3lV3p6rIb6zyCSayzrFPdFYoUbxPkoE59SJd1s1bGrLImoFDnH4YvqOgL8Kg5
9o7DjRoDj2E6Ju0n0cYTi+z5A+fxe329OyT1T0nR2OVpzTLsaOCmPwUjA5GC2oU+Tdi2E5hoAHu6
Zn2pUppjjO2+QR15TyZLY9KDHW9UAY/NwRgxJIWylOrDim/gFRn4HV9T3DYaAQxzs4lCC1KPizDt
Q8/IvppWvf0VDQEQlHQpe9zKBHI1clc8TZb+h3A4WFvht6G+1uUc/cJfi+ELmxiC9zGX3+AA2uvx
VMgKALegODLJOXTIqwm41SsMwY4m1i+V8Us/9Qcro5ZVfF/YHc4r0wNxLIfNN+KE/t/gYceSemBS
6OX45mixd+fcd6tF2znUxXcrTD8gW4px2Faiu/USLSHjHEdVDas+E24+KhdmnwitT+DcBvD/mN+i
oyK/tYv7kOnI5EJbDHvGXSPc+DhSx3tMyJDlRpAdeP3aOP5BQpFDkWLBvy7P1V7wsFvl9lCRrbeB
o7ESkMUbLV6BJRmiWXDrvY9+0kuE8RCVCrh0LV6AEVzvRShuFDXbhP/mKpO3KYJDW93RXo2pA2nv
bEcj925rbw3iZfoojG0Tm6vo7kmVSL2A4/K4C4jI9MlOBZ9+n2+iPW5SIDaOnQBWPYJ3KupwH+ia
/uIMCYlXU8UMlajoD2iYljClYr6HSqGeowlbfiO+UHdl6RJkon98RzmocFaJzcxXfbT07HvEd0vW
tZ7myGSt15m95vueRcZSPFtt4gTCTU//Q/i8kNUa3KTPoIOlnt7qRHYz8dxv5EUwlOTgX+EX6jNU
9QYPtiwNaomwC8fHBDacJwJBQ0W073XxKqdrEelGNBrgmLqUQkED84ojaaHXg2irDDPAwXbvb1Hb
imN0WiM3rxFddDSlbhR7i4P1uyYUx3rRt8TIvFkwQYqtYrzBXY5v6cjC6Kua5jCwX4C5c2RO5CgQ
ZZW89hZba8y7JUwP0LddeTOi4NEtObhFimSjXBW6D2st1b+CixwYbQUaPs8anfm/Hn089jPuaz7m
inXei4riTD5DkT7U6bH5IoTCGAxC/pB8eXxtuDmvHxl6MQ4oEWX2QMxQA+ygvx/UUEZ+e7jlZ8MJ
SI+S4ZG7FKq1QjjW2IWbK4M/FaJwkbx88rmiziZiPdMRLkzzU+86Pw4WrEj3qfER3H3AFxRgsZv4
UXhgTDezfjd2+lEwrcLfBS0UI7gZW9qFHqfT+xV86GUumf/zY55SaDZUGxa4YlLiZSv1A5BGN25b
7A6ZXMVih8tNnblNNq5hwCoKw07ZF/nxu5ZU9z74n34xke5BvnAqHd1BGEJ8TEE2GHHNWFKMZJtv
TlNYQTWVqorvhEtUw1fpPshUuAAPVkYfrSa5ZAYSweuktAettvrFs68FqA0YLKsCOcjEEwblLZDh
ByzJPNRp8GFWDQdMmid7jz3EruVKBPkE8kcdNPN3DSqa8t6z41Q0yIhQqu6RL+SA0JLyTj13Jz22
iLnnldAxmijn1AxVmIsMivJuSfiGHGZikW0uNVU6bOyDPOHOvBqs/qLiBjeFKATBM8fpL8eu4dxe
mnZeLbnrxBpwfms8IUX74Ao9KrjDQ362jQlXuZEZhcDouhBI0k/9PrghBXDfAcB2TwPTckqx2fi8
ZktcbVEaXRTwFO2ptiQq4EMETv/hS7jql0igEwwqTCw9CX4hNglF6R86qrr+uuShIzIhqdxqvYsF
qdjkPYHB3fmTl590WXJUIYgBdXJJk77V+SNUc2EJubYkkdEo16Go4kTBh96P4qrChPGOqHPklRUo
30vFAFntcK8iHhG6i6ZXYyoT2Fco4pkiO2Uv/Nell2XilBaKff4gpVeagYD1ToabPDhoXwcwwPEW
tdr9ZgMhKnKUWqfstR5fzluexDdj22thRMYp1xmZVNoJq+lZ3hmQGlx9QvrJl138GMvDCSNcBvIh
kO44FJ78hs5AeaAoVfnBHtZFhfZvyvrw7hv0BEeeu7Kv2UfaP8uigXSCHQ9s2cSFp78UAkzgjV4b
ogDVYdMTWhlssXPRiLddGErgJHSy82cKVQYsNU5az7j+NlrjSG4/rH6n7JuMoKxC+mpt25Vht5US
Gngml+mnfceJ25OjcvWPzFOV1SDT/nWSKT+fC1oigU98GWvKGNP69PhW5zz00gCgY7uJUbLHi1ld
rIavbN2TVU9Z+KuTTgSjGupqqC87z+3GdURRsFwsAGHMVppduukcf6daYeBVhwV+yQtKUqDyr/8B
GAiXojNFT4dpIvNCpdlVWFOA3Whb/LYe8gmUG2elnF1DPWvyuXYFmr3t2N3+if0OUaUS3wwhE1C3
NvJHhiE61FKeHcvhwskiJfsSeABIw18JkyQjDHgBuiBK2fiv6wttlzBr8oyO5AY+7PmnxmLqeNnn
iZcnO9nvRg7i7koXbfmerm+eSxxbNF84yvHlV0qwhE9kFWOG8wkp+TxBeEMONjbm3743Y6XSeRQZ
DsF6vgivgnNEB2tFGka6eexDJgD57B5fjKTE6TUw9NUCd90zSuwgdBNiEE2ffXgxT2Si7FHwsTvr
VkCoH2uBm5HRa3aMGcm4EP2wZBx/lPZ/6DG48g5AvjRTeA7T30MTEM7t+P/WyW2iqmrGOuErJb8x
coPMREUBCCeuepiBLl3p8DChqLIIsIrFOnfdBE6wecr1xIibQque57G28fVHQlRzWTTxG/TCrbkJ
M294YyaWlmvBxf4KUu+ifKXjQ1CryXdMYRFzIWWNm/EEiPBVb6to5GoP8SfJJWL4saV2+xCn044I
ykYAyHlwtxfsF2Bqg7YcrhwQESHsk+dGncKILAk+OH7wIakEv6Drv4BXwP7WVZNc/SsGi0zcxAla
ZqbErS7I0DhH1NRCnjqE6coq2xd5jkTYQoHgt+P1g+KisGy1r5aPJMTrQJ9q0qAYjNCj4LI9MfBm
gELXl4evI5bUlHhD3htv8yforeKWvhE6MqGJ6W5dUkkES40yT/zFzeL60VNd1BZUNlJ399aM/gA4
7hnYPZzy/i/AjHxYY5yv5kRkNk+6mzYUtyr+df+AVV97Kae6KR7prEc3MiL0xbcX6PY6K0rtXay3
KlyNmEwXWBMJU5JgSWwgd/91FKetvdpEqXF8jNqkAStkux3/glqjpw90lW5DnIGnPtCI1bsPhxfR
Vsre9hTg4O4waCrnWF/l9zLBYKSPVpAVbQFqzPDgOqSorFdlNg5Bzz6TkFKPQmNFx44pMRJxI4ag
Dor8i2ovyOaFkoRgTokIKe7fr1iqRwxDET0ZoA18muBRyA/H1b3acb6kPxB1NjK3L7TJqqBem+jR
MoSL3KwC9I8XiazNNPd+0JG5hQEHNSl1Pwf73i1LQsUu+Fk8TLPuR+2vs61h8FfPWGG4kxmvWkH9
LwoXXvrH/ArnjKMDiEZqs6E0qNFGibeALP/LypRWvgRAZdSEtJDAeHdV71VfDQTjhjuRpQcObS4m
Qlrls7LCMTS4PXwG2nW0u2OJWbhSjiBx5ld3Myy+1FhuJ1ZS/YDdjT9OhtSie+U4Ojp0OUfhnClf
xITHpQ0H6J5BYZcfMVGhBWxKt3pWN8HFfBf4VHLQkKjBmbmqmRG3ECsRLip9dOADbt9Fhwuc3Eax
F+zWrDCKitB2eea4C7Vp0001IL7KrJBE0NwzOtflJ3P2e5JY+fqm/+ozzimNH2xRz+VDch82Z+3M
ng8m8U/FJO8uMpI2XMLta+XOi/bJDrgNh8KdrbBxE2UkRY78sETalGzs93Qgmg7YM8BQeRYn1epr
31kkAYc+FW2WlRuvUsOl9cu/ZZGpZ4cjceQbxBQxFOC44m8teuD5GTr30InYvEJGgWqkXcN3FJF1
/w6GqLAbt6uVdDCo9S93TolcXSjH7wM2wbp8yjfC0hlAmUCVCarHwKqAQlJ/EP0PIcokyTNFrGtn
ZgUOkBmPXv4jHzsf6oVqKpu2QUKChccZUdWemDI9rX7i2VLU0WuVnPEqkRUBqVInwTc6mWOTVPUv
oRARZzzucRRA5Zy7Xrqh6hLrslLuPphNf+jtGWWr9zy/kZaq7FuPSa6YANPkKDkM6pGktkXcoKaH
5v8ieeCJSKgiwZ73sonXJ3fnq8zmjUJKS+zZUlZ/vnoa8Dt5UN/duV5Z+tEzUIdO7xHhioFDYowN
mOUciVbYo7WsdcbGmpsdWJyzFX+BEaj7OEHguAnw4kacLKdSwhhu7ixX5hh2IupaB3NZLa85pIf6
455kqfkbTeP0HwHsLQFZHgkNkmmfbwJHp0aMBMdekDNK368QFnlar46nDwaKe16EvFVMs+xE7gIh
RC6xOcwXBbx4yaP3xaWwLDmw1NK0R6lgzAxiqb41I6PWJJpUZsQCGD7pBA2uQYpPcAOdHN7lA1aY
+Dwh9yuHaFKIL0CU/ZnU3m1Tpg5fbW6W2E+YuxKc1v8nO1KCykD9kjmQimggjDXve/BOUgi3io5e
ajwvFTrg3eiZ80foPdS0LCQ718lPGziaAu1NY16brExVsjhqwskdMF0LdtUdYONTSlbvUuwg14hi
igzi6uCXbaeyVPuF6QZUSVDZS0iUIj4v74OBcuVPZkHWwBvCKNpbxy0HCK5bwoCJsyaHV0f+gz4W
qy9BO8oXrOoWz0xlRE3TYzDiFaL22dV6VHt/UKSlLmPqOVjbW4ouQaWCsiYJW76BdgYF/qjnP20e
QKJfupRkppRqoBaCAlGO1P5X0RhDIccqXvRg7HMx9HdXRNCqenhiLhcoqmJSTZL4TAVzFfq1rcsw
S6E1z/Hpyf3fxWWGUDDUE8wKX1tdd1WgMHjEphTddwRt0z39bKIVRD+eFTRSjJ5X0Dc5IMqHfEWp
VNVPtGhB7har4KGzDeBV53qgebFm+HQOvAG2u73HFTBTAp18iswyZ5Q2UQz6Z+4arbNVcL+zutK/
2BziKASPAXOOn4jUDG4G6RWLesQ+AeAaX2WzBgJTM3pWAg98IyXh/BaEbbxnf4Ie9hvuyvgn5amV
2UfTsxXQ2INBWxnZHpIJ6zcxY3KvK1FPv6LUIOaQhe2nL+5H1n31Tlzl6/NajnCsxafRR0OQCHR1
wjsV98buRsgCV/hWBn+OQeL+oZh7XRzSUJNsfrVZL0EA6tNdp6F69XZHiNfdYoj0sUUz8QtFLraI
8N6X599FpokMXkQYM7xl3aFjWee6nRxqzSS86R8MXRZCGe8hFaaq4pKFZYHcRtUcDrDy4Ca+5Yi1
uyr1rKxO6Az/tUsH6q+PsAZPcEzK2UrMAtQ7yQAZSfLSMhoRnL8TVnHx2rVcwoXurSJa1HaQDaJ3
cbhWntj7r8QwQ0tXTsI45ILQnc1OrkofyEcDqxgBHV/I4LgwiX/0njV6iK6RXnzl6LfVqaEoIwos
DrLdSkB3UFILihXnh0nW0njlN9CdJh9SUnx7hL8UHTOtmeIG6mX5kNTa4eKXVHPUS6OCzYX52yYV
jGyzSL1VkuaHLSFyyfDWvnzUg4WQzy4Kg22E0DQ/Z7nQk1rQhPq0ILdAub30xWwKU6QOvLGmr5yS
zd6ACdnsSrzP40keQmpM8xQ56+NCYqBFiijIgBJAety7mNYOZ606buE8O9h5vDI3NF0vddaeg/nh
9d/2IMQH1Y2dLhjQCkcEQTgRm0vRABWl5Z9u41uOhZY67BBpFrTP//U0Gjp0fWESEHQQtNbH568x
KjIEagg5Hi4UfnWzIAun+52gt/Zib9CFr0bIUS5Y0YaVuZLTkBDaVW/lWXm9AmmO3ZKw1MBU8dZu
ClMvWFnPIZ9ruJyQs1Bi7QYG4AYIVefXDimGq9FFzoPhCn4nWqOHisuHibAy5ZdQ0VM1tVvhodTb
22Op6fqJxC3JF4mx3RtA1e5WfkWoXjs1ME2aE6xrxOpDjwVzqSUN6/Y0lxJ7AfkONigxDoBDZ9/+
awH9XZdWPdfFfZ9hOYkj36OOEQJ3tZXhOHXgen2mDp1j+6R0+zDzUhi8pwVAy5At0rFseYEbJGde
LrO+pdMQ+Q8ywC3VNvkwOdJIq9/1yOgeeTlHz2V7cGCUqkwVPAsUTRlbPp9yIP/XUloJvUw7WdCo
1Utrfte5kTb4qFSduSCvc30LxLe0SQOOTxxmjgtJmjn+JcYuShzwU+7MFYMROjJ1BGy9sZnrQ65Y
2YeqeDqFpgR8BVRL6+7kpeJUh6XlbuOEh8uRDy0bNGB2nPx+eUePi1EMGjRna7LUCVU/uCQD/fIl
DP3Vj0DRCxSmynEocUK4trWXnusmlnlrNe9rQI/gJcQpmwRUl9wPvC6tH8vfCFE4yr13GnWq+KlL
+Rx+/SZDWmShBtYhQP9rvpvBtYz1V6QlNCPD6ZmGxYQSXczUqGPCmUudV3rcaRarziBIIsF4dtoi
dIgnvY5BF9XITT6keJKejilffkio8M1eoJaUkuGTz7OuMalGLTb+Gdc6FqF6ASzLHaZKHXAdYuc6
s17p2IeO+5ek3Q16N5yd81YG4Llh17sbw0OTkQ1PV5/ke4wXVE1n9GOqK++EnOX1LkvoJXkRbpJ6
BvwZDQgGzPccszugdSlhMeO3IXHG7+dxVqMSNz4a6RIsLoltnSh2aHjDXMG5uIMeyBkn4qdTpNK0
R2F1H3bx0yxYRZHZvxVyQJqfcPQ0wUMbGesXz+GrzTVNsaJFg1PtDSEp3fu4sEJmQ+jqM1ut17qv
rG+saS/rQ4JgUSfw3bn5PSDn/jw0dmGJXeKjayu2yRaYAz4SYLteUkDfll530BSz21eCWrnSshxJ
8I6HgigeedEdIP5e6tT2qboPI9/G0fCGN0wWJX6yiPfqrwB6O3sXbbEcXZwKPFQcre9Y4w0W65Gv
Pktilg8VJ+uAly2tJNsjiSCeeblHMSCuFzRX+hjXd80SX8OOL+uqcn9RxhzjgA7TbOKATKhkjX/e
m+vImp4GBVb0oUImu8GdI9j9XHfrdI6vRUk8fMT4a97EnwtKc7OwfgXnrRHZ2mu+dV0jZP6IEnBT
WLOZoyzyixRxaYwvZ7Hp2P9vC6MVNpj+glmgb5yFVOewcRrzn9ydDOXQCHpOzdTuR6c6NaXXND9V
WC/XmU2DFS+BjHi54vPJI+uMZ0L2gLhZZ30gEozhOItVrF/V7elkaOjD3rqesRtf8qeHhb6eIum1
WmCJBIyO8br0hREf3G7RtRjFnatg4Jfx6jI9bfS+5oy6Xq8OTnCvJokkHc0oAP8Hl+sNFrhW1w3P
zj7olRMRBpg5TIoueAB5BX856rpgk5t2Q11Q4FIY9ozlx9WcbitQY5JaHYlIL7QAL6vLVM4TvSDw
c6HDfpu0utxrWAtB7MmpSB7bT7JyQfGhQA24fO+hUlFMil3oX1jloOU8oZoFm7jwqfOUMMhjeqNM
2YFuzWh0zV3xhVW028DQbLlQ0rK6aF0VNkpPp3ewWp/pJ9dNmEoKbwV7+yRKgFkb6seM4AfG66qw
AKwU+5r0gppVWzfwZAMYovEw6V4lWSRabzf4PDDSfvYGynr9f7Pzw/fiOzMYm9DgbIY8AJtGF6Nc
+4JfksRnQg+UUEk8MHI5lxX3ZfGSWQ5X8Mw+wV/QmnLXwAmgIIKL4k8qq2E/Iwb9BLCmS1Knbna8
Je0O6JSKf4uOrpfa1lwX7WLefKjFsCwVF66aqMeGhj6gA3QhHRv8t8w9l0fmKtIi2wlQyGUYZyNZ
6XytspSIr7IhuoHHiL8lZO0RvFDxNoBdDFF2a+GE/ncrSMtmD+LNv6rxzs/2VsEynViWBL8qkhym
pcVnlI5VNR01U4CEeBKxQ90t+qpTTyG8ADE9swc3HhUQHhYWZO9yfQRoQ7DA+tgMt+ERhLljTY3X
e2/ltJ2SuB83l6qNqsRmmnRNFNozNjuZwzk7/jJaCjGP7Iz3+eUICBHdECI8zOZXqT3jg5a+FZC6
/Vq4q0F0O0PZhLlwdLbm6k985GGRbj4O1XYsuuD062nZzZMJianT4lnb8K2qXrcE/PgWshTrat5k
PsrwR81ezHpM8PFLAEMIGIBO4DZBdw3TZNsNoicAb0xq41UpvKHAfKI+6TuA2tCBtg0qrRZ9Z5Xd
1nj/wRkdwmY+WQ+B9tbU4x4LAXEeGZMMXl8Rcrbu+F5Houd2Lkw4LxeUZbsfcrkVsRli+b3YfZC7
QfV9dxeGoJyqimukYX4+FGiyBcsBVhpDYVocwUwGzrmXDJIp2h0AC/xr7numm0oxGX+UaoD693Ab
nsYKK3905lj+jLNN91UUP4vqInZlPsBrNo9BiO1jj9t/4IZfvB1IQa+8PZLZmtA+/qQjEDERBQmC
EOAhrvq8hfg8qcWGxPqd6IS5Ldh27GhS309z225iMiMCRQ+EW29UIx4nYZ/IRpSiVFXiZR2ROZUK
P+FMBTIKn/I9yUd3xvoE37wZxmzhrro/ZGRTCNtshLcpqBl5oNWybEWVte9T5H9uqOkE2jocKdHd
zGKE2z+Lc9NYRYut8NqlPUEO0AiwGzp3OsXyawkA3BgkduPIl0JaWmDWY6G+RJ06TbpoPvR62V8a
j1nOMxjQNzJ/Uz37Hh52O6dAiYQXqTecOUp0V5o8xpHO1bKBzq2vgbXqdDcaXXc+vMKjwYPpMzfm
vfcIgDJRJeMCIps76YgAkBfymbJJj7N12ADAngqkxmHeuMCuc9krUdK46aep0tRDD1lw4Xf5f2VG
fm967MT11PUINuVM8vQKI5pqUohlWJn6wxu6qDsxYQam7Qu1SCv7plfbJWYc0juKGa5tCCcaq2g/
e2Pi+/BQU7YdYfikWgn3TUBTXdDWHQOkYoO5AITbda9WPeSncdZcrEN0lZwsebco1XMktuFmcba5
wJ23LeYQDw2PH+dqtSGC1c3RYuggej+f44edcxW/7ioiVtSlxD21xU07DFs5obnPC73wQQX8JCFW
uvJm3+M4S+Gqpw38l9oQ/v4I0ySbgN5F+53tdnw5BtRhOxduuXl8+8H94nzwQnxhypd7ZzZtSr+7
mtMzZVNMx7cmAPeNwoI9rVwFRXal8G6YIzw0ZHGDcZB5SVceD6K9FjBmHmP8wupU1/Cff1Vd3KYB
XAKTYa+sJfUq3aEoePwMrjxJ/jcxo0Vjh9wcH2pjCmcQku99PDG0fHaWe7iwJR4j+Wv3B+L+9jcJ
EpjJL4fgnCgDXrJSXeWZiFLIVvMn50QLumZxMu/x+PtdALWGIYNPzsLqsvZmwdTkIkhtpVDT0TWy
NtAP/+S8tLBMf+a5JGfJ1DDL/QkyGCfrZnuTbSC+Oa2r/mu1qhlsMh1SiVF+pzhx0yTRS8PmRbIK
R0kwZpryh2HvhWHytMUgiMVC11tzdpQWn+1R9JYHcdvkwTNNLoGh0GA4+aepgnTBGQSaBahtYZOb
sTHx1xi2nSyZgV+gvSpBknEIfe0QkO4CNvDr06YKvvTVBgumwo1dCN8fhd6ti5Y8kHIllgpldnMh
HbtpJiXv2aWRgqS6VjOVt5XYUj6itTr6EMNRVRwwxDggIhb4v3F40vmoFjVEIVag8pqiQN3SJmGc
3+jkaOnH4oIOtzL4+HJVTssARk62zyXf933hDUizqztFyG2GYc0uY1kpvkBBkz4pzU5NHQL0Jx7j
1sSjsjQgd/GEI2tEXOaE+hf5RPn0wsa0vGUd1VctX6K3Fomo21Emp3kc3qYhxXynZSss70NGug7K
aGQUaSaWWSHzn/dO6Y9p75CgPTQkZhVM7GlbzdZaqd6j+BWnqK//zE+aW1FOWmcdSjHC7fhi3lMw
kGr4Bs3g85rNra5RtUJ0Jjv1QdwBqPEeTtIEBEmqw+yn00fk929I+8mPt37+9fr0sP/zrokoRk/P
O7SFwm1NPv+QEeoU+Bflm7J5PIp9UCBWaKUUy1q4GnyNn0sEFJJgeVk+glWqvcbA9g6y9XLHmIMw
xmjm4Mn/no1G2vWP06bWFADisUAqkEEvlA731+EDXM6qyBVQE7IIQvkYyR0oBCx4AaE9a42iemO6
HX2xI1pWbHsWSusqA7DOuUdekTnFJf9RrA3XvfLFwlGN8HK/56v1Nym1w7tP7hfmX5HgZa1zyro+
VBXNc57b/6wXjGMS7KNTePNi0vhOunPjjeN5bNMoqAe+Ch1OHuhTCdUTZLVK163KX5HtnzlZjEvj
MOs/+MzCWPNthlD+ya/8AKcGRjUGxiEzgmuN29U8x4y3KHj7Hh7C4B3huELZpk0886+F19U/yqJN
PKuAyGwj/RxZAi+daaPuuE3lmPfJZi6w8RMzbMImK9LwRdfx5NN8x92pidu3ZGAEEHXT92DG1L3O
V+ernUDNG+Zom4Ph8eJ5zj5EVEOCntl42RCRNNufGc/zaQN75cqAhhrnikOGA/va/mbSDa3ibnHb
vvOrEUUhYL2cT1cAFwl0rxc1XNYnqcMlSKGu8+ZqfJtL9rKywc8ExL8Fh0NFmTqVWQOdD11PFCR8
P1AvlhvbtPaBa6dCToxXjnlk/kzXzrfiyqrWDGY0YsND8OWp2q3lV62XCuDNYfb+w9NQLMAFwrRX
WYtuVT7gHhExNzKgO6oOJCtCAYWsXGU/maytH21gphj1+RmSFEgbS+dJrF/5ze+OqBft0PoiFtKN
eIuDI1ws0in9Lsg3oXVqc4cpFRQuATis5fUvJJt6hwg4t9JmLUPz2o7iF2pR6lX2dp55sGF4e5RY
VBwbgQqYhbKNQIvQylHTCTlGlCGinMb7z080bv9FK8rX/mdBDzo4VMQC/t9hC9z4pgNnIGFOpr/j
RKS3p2G+E42CrJS6JeGgAA2Wn0nEeG/tZfJM3wnwUksduQsl3bwIyWgdMrQpwocfT46awo1Ro2bh
wmKCpaviUK+9IAy/6PvRZ/gnBcHR2OaptwysuZLRtO2cBRXXRUtXiNLvcjQPfS0IG4hoYc2u4oEz
z9gFnbgsPYoX+9bwXIiY8aGFhIsEpTrzLxIntoVR6KQZCwx5Po5dSc4BH0FKhsdjrezkAMZ7GzFY
yYNZh/LC3wd8xJLfBQcMlalvQloNZFVYyP83L4HJ+vSDlZRu9JFKC+hYkOu3YqNq0sloQyvHOC/0
lWBH5kOPVwnitiX/vvkuTf6hO07JPnL793SSw/RUX/AJqDT9rXgMDEyWOqOYvoDdjXGtL7G4+JC9
f8QZaXhnXNU0JeKzxohzdpJXqnhHHDaGm/HYO3mJ+9GRPxLHys23gtm0lSWzeWgVFwIsfUmpXb7L
02VAkn2rj+oLV/gdAZGWhWF5ifuAYKHVlP4p8z5py2vFeM2w1v7+d0vpT7MI+R2t23+HE1/nHo5d
18EZL3sjDEIqH6+hyPBFOIiBxRWPjUrfW83jmlmWGDp19fklheKrQd1BNmXu0S3LJTYOs2Dx1b3/
Rvy3SgWSPHLWLwNpgb1NHapUgXDJ4Qr5UfYNARAtaiaCJ0+iH3tWxX35VvAjJgOS4/0FXIiyhBx0
lw/ySYid5T/pW5EX/J83ZU5U9HG38myCfQU5logcVGPYdl9l48A0G/JTKxTOnZvQPn+DJLsWx+Dn
akFN2s3zVDmQloYbpeGGWhftVm8VAWVt/g9+0G21yrAFk+U2rkP3mKiNZ7HySK+3GywiDt4dRUr9
QxXS+P6Tl9lwyHB9IYKKDf5mOQktZI9SFSVLexUQPgeUf4iIWB7J767SypRPd2rkvrjvKh2wLqrZ
u0SS3RtFpLQppCavRnClIkmIvZA5jaBMygp/cGqg75kdx8Tu+MwgzaQPbQjD5gVTrQVetBLQjX7o
NBZUKv41dF54QxQHq4L5Fob667Iwb1t4rT4ViYlARVb6c0LZu1JcvY6qUkK3i49J58U8JqTADj5c
OBpytDeutpVlb3VOxl5aWGat1fLbUEf5m/OSBBRrbgwfmQkiFlawIJ9VRJ1C68eYpiClNW0KFBNo
l4NQNvFRy7OLg72SYe5G34LX8qiDIi7ZyBG03NU0tzynCpaG5kRgUyPBw2bhAs2lwPK8wgVUJnVS
Zqm3V3PjHc075WxgJvFc1WgxvZpa1mEz/V4CaZvHaj+47Wlvgj7Pfjg3sVMEJBuEs5aybb4UwMdw
S0Sdtu/g6WBneQe4JUfq/2jFcRF8MSlynqutZ8Uvl5zrDiLEgqqqn4/ICxfvIEUmtNt9jgZjRsiH
SiBsZWpvpyhVZVFyRqsBXZD7IRosUAKV35YgHMgJjX4Y70QoKMOOdwjJxz/uhZRpleDNlnAhuuxO
Bj8iW7l42Orbnv2+kJUDQDJMDmQTS3BJgrhmOUspqDIjZ9d7JEeaMBZK3nLB2QqEx2NIh9K+Eax6
Pkpn70QMuNtrwcx+goywi6vEDFl1M6Pbk+ZRjMQA6ZBV/YpuLrtneU/xHuTtAjkNwuYoOqdRSmZ9
1S5iVbHh3N3t2/AhRdA8Lr+WrH78+uEWlp0o8O5qhtcIW5IdkcGyzU9L9OEMd6S+TKBi8QqZcgvP
jU8tbZhbWBVBOghmpJ90VTE9yGWbk4S1E/1VDN84Y/n/pOOJ4bbkI6cc6Z26SkN/LnoAFwPFwlrK
mn7p7n4bdR1jkPFlhQQQLovNRIVko96vf50+xtzOJBCS3vAY2QoQUIPqC9B/QKIIR15YlPcryIB1
gT0bVGJskWsQToYl/chaHZaZRzG+4q1+YVioAm2FlVHt2jZ1VGv4Ce4O4QO3GmRDcVGnJnGLKS+5
E5UULPSq+G5xPrIdWXLGIXsNFaYKKTGfObR20LpbJreyW0Joh+Hrd2Y5HlV0EjEzfvTdNfQv82Sf
qY9XZJ8mVNe7KWrSxDE39IyuEsz7diHdCBlQ8GrMhy6ob80jdYeoHDyUv2VeKL6KEEP+ZVQfFTA2
xbt5fv+bkALlbMNwhayWSz+ogkZcW44zYUrLc/1wwceOl6W4fx4L0YCqHLHmL0eIPZ2PHhkqxNUX
GK2vNZ/EdqkeL/E5YMXbdwC5WoMBCHZxG1+XHlzfmlNCOgmzD+dakTzyMD1QIsEJP/Wh3IvAF6Bh
bgj+M2KXXqPjWGuaBJgP/m55NphOkRz7YwoRoIg9IvFIjOB6D92LMJg9yiYcsgIW3w6sGcop/t9t
LDv4FhJu6eOaM4Kr2g1s/nOBOivKFFCu4ct3sE01dvHhYKNMJ5L0VKKXUK5koNtZRONj0oAWtGBO
5Wp6gFxrmWdHnJCTwrM9pDvdWdUpHfL06gnGjt0/cV1xiNy1xdiYG/f98UOoe2Y6NUD7ePbOktf+
LQiBzMkoFPQKP/eq3nPqQnRXcYb7TJLc2cKuSFkL92u08oGC1d6L2A3u68e+Qc2o8fAXj6pnaPVV
BWkDRGXCRD+drr2bT8NK0urpeuxxtxL4FKakkanjKbe4EEgerONHZUpohjfVFfApvjpJHlhjKxC1
Z94VvxSQ0oqgID4ngUS3WRZqMCX1wuzuTOpP4/s8KDnegElBSN+UTiA5faI4J5s2zerN6nCVPHbS
de11Gy/1LXWY3SkhDj2QoyoDJc7hU1PDLVGyjkqOlsFvfIZoNd5ka4eSvULFSTMo3xT/9AgPN1cm
2gxq6AyJoQokKjo6ji2qlp9PpVlTULPg8hG9Ei+9JCcLkk7lweMGbu5y0uG6+QRWtnk+SupGkRxK
SC5k2fOMiErw7h0CKn9FZncZH61z+yTS31hwJsHYDr0dnWgNxumgwbE8goe1bBnnjdd+wCOnXdBt
Fg/ZW4JvKZL8tkvLFdzK5xuHS3SVSVj1KZwBSQG0n4ILwj0CHHu1z4lVmkyhgtLzr/JTlllFj+of
TwDt5VzFJj1c3RXUgIsj9bUNk8a7i3yFaNZiEMEkIlE5cb9Jw7IkQEIwuC8XOySaFZ1pddc++pWP
MvFEZeY10WUezw+8CVK9Fk9UMvwb8FGbqUo2EWA4LFXj/uHkpBrnlIYrocyWRAQC4nzpDQToDKmA
0CJ+glZ5ZF5DI+6t2nCoFkJ2G08VOinHSWmYHrQoVmTUqbc9jUb4C/DeRfKwYyKja5fXckQ7koSR
Rp9iQn3IFWM3LnXeCZz49tRbGQLHpMAJzfHb3wm2f8TbO1Lippqy1YpfsrYXgi6hx7wFPogDZ/CS
X6ObCxXsACfvGOM5s9mCjGRAyMKlpcj9/gPhTsHC8jkZQ+/WT5cA65MfmlzdjsnkvS6Za3i2tAnB
CdK6Oi3hn8pIVpvBT7xbVESIrzpzSWgYWYFgQgqHrLMqRC6G5W2/WmmnKuX2lOuNWXTPm1dA+xb6
qvkEpwImUbVhPr8c2zOOxYP1wblHtDgJRQGI69wP5i45d9NK1HVZIg22QXq3GwtZOPv6+9145iv4
KSuokL/0HaQCb4vfzNqS/Aq5paUQQn7sF+NA98JWLRts953cWQ+AkT8N6JvLQ4MZvydi5qIIi9+/
lb+KP+ntd+y5e8KO3sNa9OuErqnMVCBi9/AzEE/ka8hcdEPjQTcEMWE/RSpHcuIkc31Fkf9b18yd
kzRSB+KY9UF3YkhLHJMBUN1fR5qtR0F1iIG9Q0OuaG+cXc2D0rewANr9m7Z3BiWgo0hbywt8qUtx
vWegH8vEPlei+9EXX0M7l8ky45txVyliHvcDrZwZeWaNbWDSMpN8xtd0kX+CWSHyU2RNbj1IjqVE
ro0CtsqTS+d53c7NMkRi6m3u8YS+zqrxZPjlF0+Ckwx7PDkrNN0CATEe8IiNtf0Thi4toCZJ3w3q
EI59hoBOU8OYfNYBli0CsFBgk1gAcnLFnEfpmwOqoFEimS6lNd8gDct9wauhXUjjaB6convQRK7k
x3K+B5+taf7JLJuYsuRzU5oRRIF2hjQhIuZ3GLFxFIhRPgBlHFLTGeDNKJ0KbKWmGzEVJEto/j+1
FqE1EzY8/mb8IYnbkODccDodvWhSyrF6nzl4263M1m5TWXoujYreWGhK6bMdDyoLI4CtNOhGnoDE
ymtZfleqFDC1kRxvblZA4wSQHSby1zSq2WmxMmTKZa/fvJ9PxABrNjMmoAA2IJINr8CB4qr9NcDp
yUUpkZXUlWgNeFnAKCPYZrAg1e7nN1BD8Anjhn0ZhPNa6H9pLXOzwtkJB/Kt2e2/Iy6yarA307GH
T6sOVNrQsAHaopULMZ2CFX21R+tiv3txaJeExd1BIi3Rc9H+xLvIEtUf1NcI19cIdj2YEAeQ1z9D
+RPkq64IxtVoOdgSXkecG526nmF+5Ct6hRnNgsGVlyKgrdMdidirgj1snouY398lzuAqZmCEuVaR
fOf9wJ7NnW2GDRA7hLv1B+5o7Gu0YLTlHj5RexAhSB0ck80WuROPrnbB49Q40tTGH8+4V1GasG30
Y0YLvPCePJWpYawZttEr3aXHe4pbeHjmdoyl0rcd+WLExD39yCQUS4yjDANKWmhd/8HerPN/AULp
ih5WJrg/R/K+VCPCVZYFphCC9sktcoITD+NjD1qcj8BWL95jcDKtpY35CPwUVYvW/CK6aSQ9V2BO
Dc/d+dsqQ2v3yPOR+6IkWekfLJo/9JEryqsVlbpiz0gy4eXG8ge1YiEkQgE1isiBsnI455Tflg+B
Q/Vk7d+LNEW0X2aMsJZVGnixBOskFqn0mPh6IxePG4+EOebg354UK4XHV2CzjukUEoAeKYKMUdCq
xsMqzfkzb4XXR28U4UlJEI4P6JYT9zYO/SWXm44zoknXz7Xyw9t2a0EnjMwBVwGyonRQ5Qrdh0aS
QXa8ll54DPfsrUR6Eo30zJIOgwfJwT2fCq73Q4EylIXlOjwXknq/Y3Sp+CqQghBU2vf12oU4d3KI
SByQNtB4/+DmvNB96r2dr66mcCjE9nNmT4XawOYKuTiRfPl/1aAVTlp+ZDqcvjGn/VxAS5b95q7d
rGYEGQt3ESxuPhgrF2N8J95delQJu9xkpsQCxMxN6KOKU3nxRzOlaItB9Bm+mw+PrXkAqOUzv367
NrsxU3l9uKuWP+tQqfmXjRNa+D3aSzMibQPsPwEsnXhwdT1Ylq9YGOwFLKYmAQlHZtLjv5ZlePDs
l8PKpp6qaen7VS2ocJxLMYDXflURCoK9p6gn2HefpC9LwENqf47Gw9G4gUMESKoIR6Af+5dxc1L5
uxVYmy2FKdQUBLFKwKa3cfT/lO3laQNJeD4PQ4ng0o9PPReoV2SRej0XRQ1RI0Ul3nUBnDKigHOe
8uVJYv1sUh8eyuajTrPyMNNISQ0xUyh/mWlBO5XvpQEdom5snFKYz0pKQcq2tyM8l8qhXy3buGHG
i/RtQ3WtCdvX7j0XiRjjHpHD6XW+PNnefai9HD/JUMdUrBhkQfS6/CcM1NO62ONqe+DbscKdUn8+
UX9q0B9tJp/taB3Q8dPPPrkKDTUyYRZH69TZ8hmGcaDGdyoyjGUW81SRX8fBKkTngKdGy1xbP51h
IlFzonyGAnzUYemQXlb2D3Bgz4txgXJl4LqhGMtJSMStn2vm7+bsSI8BhOG89ZmH9OuoT+nYT9te
xvwUklqxSHF46wQy5GOt4BDFmo7+hb/8ryctEyoxFrzuoYrcsXLwMpB2pHn1coE+yLA7GknG8wEq
bgLe3EEhVWaKcRZLkTMqS/kXgOarUq2OGAsXeBTfpy/wBWlHxJ8wd/ja9D/0W9bQj2S14GrZccBF
J2GdG1689D3dod0US6NILGLIu5g3IJfSj0poVwxfUdaighfihj/KL9pidEzmFIU1UGruZ2r4nVFM
uLenxZwP8iMCBmEiQXg7qIC1y/qyNZsjdrlR7h9r3gxoiMFQCCTeQvhKVQ5rsCCQHZtuQ7ZhLpNf
qLR2Mg3plaZBSA+nkOXlSy6UVwetKZpO3DOsV3DW+vuDr4NZhsM8alQfFym++uauFucBViLqhFPw
9N5wv4ZQReqcezMfAX/l4WGVaFD7EkdTN7eruWdQzZ+/oiu0uSuF0+8SBurhdoykEQHdCXm/5WZH
e5DvC1euQlv2GXhg2exYDyYgLJKjazOAXHez3eCfGkXV/CJA9biIht60o9fHxDpqM0d9wC3zsjZq
jL8w8HAztY424gIIP5AOS9LMSaPKvJhM0ggmdOkywi+jtJ+gPbtt6Eh9VeARQtfkJ5YLsEtqv5LH
cI6AMtZ2ZR84xDba4oz3Fj0DO0/G+qT7fYGJpvpEf4kPqDubvlbH7qHf0U13RR4ExzSSheO14Sbl
160II9mQ82wTZbzw7dsPh3u7ceKlzoIL1SaSln28IQqpkeh1az0ZctML6G/NEc7Ycxa+WqkBsFr5
HGB3BhOFCVqQ5gigcA5PriBLV8JU8O+4U1RoihaxOhUpEum5bGZOXre9ModkFDY0/Qqq2H5FKgeq
U1IlKSjLLlZP3ilIzAItEoWl+x5DrEEoKSnOtBtWznrO6qtzQPYh/eJ464/IhTFfhP8jSR6S46eX
LvaxG+mTruLj2CSNMvQ6FocTDAFqokrqvnro/c0ve45SBn3UoW2mSi3zmEoJPUvV76nvovn5/9zv
y1IRkT/nEtn1A8owULuc9u6Ejk2HXXRUj8xZDmZbg2o9k8vDkQ9fjqL6m16I/HE7Xbt8f/TSXnHc
gQftw+bi1c0YlkQ94B39oB6IaXfxxxL+jeMNT+QHhuTv0b1Vxw/JEJyw9HSGd0HGoXp/RppUxPKI
ijMsl3RA4twJdadZcbUb4IZOID0oeC/pSh/7bsTFgIMw+Nk8FXUU0lkCWC8h0g4OBn2FqZxvrXJt
AhGfa4Cp/fLHZzrJcz9MVyVUEyfyiQQB42Bk1trygy4Wv9cM/bhUoIjvf1UqF5W/p3pt74ZLvJxS
lSQmTHxOyS49H8F1opOo3BSMBWQPBoqR4zoALX7IXV9Q9VU08TxvDBQXDcpUqeVGPcqRgzsaczre
cx8FZN9+Ndrr8Ec0vQO9Y6j4dH2vgp0pF27UCmhqeOvEajB/Mn17B+Bt8ORJnokxW1p83QovmFMa
fqo04xeAwCRSHUhg7CVWquQy31TkFqc5yN7+R3GFgon3fLHVU+zbpNNDgZ5f/i9bI4h5XbHzA441
GoA8ZTNCRBc78wEfeuOkEuKKNRqaJlb3DsH/lD9sElt5bmWuxfdzRdsW90+0mVCcH1bOvJfKwJPb
zCn0ku3LHwAotJwP/ImwsvIP7SKA8/81XPsBm5eZnRKC7CU+heWJv7KAgyHxIQ9x3abYZiA03Inj
tNwPGACsoOkRKckio8D6RGM1lfPXxwxGUej5ju4k8kl5NZgiqGzUnPtDAOVQpgSWGhgIHy1ZpeuU
ybq8nWepu67KGH9OJ/bvPHrkEOaCIe1P4eKvEX7wn3DAbT0jzGMMv0UTdEUIO2wOJ9Bej7NDP+ft
vo3mhdAi7J4clXZUimWXFOE4qGZ3ySfntZObHfe8IY/Tu1ejA7ft036lft/aIzjDW00NGDSjBamk
1JbgYKfC6VNk+KA5pexlTBuZ32ouBk+qFxUgyKd88iiw8imprQ1s/iFg9CJ4JuoKXsyGYoyp2W1g
2EW+KVprejIAClNIO4qL//67X3H0InwtHu7qR5CKGiw4zmggYTPZTiZ+5xeX+7lj7yDUlEJvNTTA
aCfpJvlY7bPr9q8uO6IbhhuvC3uK0yea8IWsCVT/1b4tgcy2eWLwop2BYi+2bJHoF/K6Z3OoHcfE
DXo+rpgCRQPYi1sj7314CqZjihvEKLA3myS4LOh2/luMemsHeBjLtGEnij4b0AzNHJT4RQ2DpErf
0TQZ+J8Ja9C8+Io3J9NbM8VcNuC3aVzn6lh9onaM+0MCHu2vZgenlyydO0vnvr8vPtol1RK3E3Pt
mW6lh6g72p8S1pCLLtN1xCJvqMd/z/xouYHTZw103JnjrPy2B4GYNzGKU7Rsd0TTBaGsbll2zsOR
QiBYsKB1LuX7JENZuusfSnbBPOdi7rRYhkonQv7ztED9ISvRue81Y5W1NfSWyERqpWq8SFEvXqro
P3TuKQc/n9NnayHX9OcASMiPsjiQblfAE074Zwxb/hnknzJrI5EnrNWjmZRiaXKTbaRqYfWp6/mC
Jp8CsBsP865hw66+EOOgv6Y1Qz+mJK14E20YJaxw9wyqddTH4j6uL/O7LS4OSqDon7fURBZkMPP/
UhL6KejSGWGCsmw75XOdM9dGZ6eUiPMj7c/okoRs+ACzuyyn1U3HTPLLJ+oCX88yW7TwJmVUp472
TSDu+WXx1jnPePMwOVlrmLhcRbk5oUR0va4qFlm4udPvrEtZ/GHBvSkDZ1KtLjBuysDMqa7oBjyh
/ZIDD8xnjukdEdzhYFHyPnHPExADsCed1YKiawSNj8RdFMT6Cu1RYhdW6al4S/t3h6iBx7ZDmHtI
YGjgYwWKrzW5Pnh0UVbqO29hweUXCkMNvtpdk2HaWPt7I4hfz/2NfvP5IEcuQgNJ2TXzNtdgmtcK
gdW196EYgnlVtN1sqpDPJ02L27FzWZA2lvSzfkF0yMBmuI0apLfTPNsLYF9lQtfirmRCdTbk6hs5
Yz0MciFEn3wCuiJTA4Stcm0wLAuOKnWo3Wi3KFwcnZW62+hvoPVJXcCVG2ddTHAM+CcfpuvEnirD
KtpCs6HOyOXEv1W6ntt4EiHvIkUqWmZCW0Hmb/seY+urB+2W0xKlD2onFZvC54YwS8u2z2ABZsF7
rVydZDS3jXpuQ79oWD0r/qzCRvqlqvsQUQC5y+cnC9ZdEdrD2B7vK/mH8MQq9dOx37iHhUJ/IT5x
WxkrN1lEImyPlA1kaGLMq5ie9eq9p2smEZg8YwA46/JZC6g0sNA5KulcMGqQz/Vm9GsqM80VOZlG
V7BqFedm6SAUauO6mIBsT7bE3OfpHsPenQq6/hqGn820yYT7WRkUvl9xadVRz9mYFYOdVPFEoO1Q
Nu1ZqBPUx6zz1BnbqlNRy5czPMMma6+aIyErZxWV4793kiL68BR4beRKMThYTi/g9mHDV3mcDB9S
NgR8oWvt+FlQ3K/imAospDRZ7BEKyvG9sK4IxD9VQqX03qIw4e2U21IPPPfKca2eTNnGot082E7X
uAwWwrGh3KJHUquBf3S8f51nJnlo5MNqlIoLeOdur9mTQHUtPsUBnMNyf50QOMwIIMUOdIhKNojG
Bo5yTDl58PGmFl5D4OltnWYiUiGbicXl4/lODf30hGl+3C43th+sYm8WAEzuXKVsFR2oXA7hThpy
AQV+QPTI/ZfsyyCvL6jyXhOA9MfJEnAkl5yHibprYEeg40yZkN38rU5s+fCd1z3XpnOqlboyBAnm
ouWS1+Ws8nSGR1w4Yowcuc8XQkQLZQ45q5nP9w0vSjGZoUCjhv6hITu/FlnUJmD0yX8CyymWkTH+
zk92AGHcwqukAgc5pTaHNzflx/QDMTFbvVm6R5gp4uy82jJxv7yA5I05E7Yo0MEqqUKp8OfJL+H2
HlPQ7EgwvzQQ9QRlWK6CMOhFwp32aODbk85WJxyR1kF3WXFRO4PBTsBLumF+qBtcS3iBlEAPrk1Z
P2SUAvFfGv3CuWuu5my31KPFyDxgQyc8Yvg5ttwAaQy04q2Q3TAYxARE3V8dacy09jbg9PZ0s9ax
CHlkyn2qhtqZ7LLE4zJtijAjSORVnJmE3C2H0cKXmlh2xciS9Dl6JHFzzfGGnsvda8WYxN4zGIK+
06DA7hZhhZvDpudJUXJ9mOiX0WIlumtO8RXp9i81sKH6GI/Q24xB4zWg5q6vuD18GJu1gEdU/rTM
cM3Pd2DC4Eq88GgbPN/Flj13jfL3wybULc/7qK3OEMYeti/27GUocDIh89IK1qkKZW88zAHE8xsj
VfZ7zOGVhjD6xiU40rcdsWrKf2H2h2ZFvNTFSjnJq9vhedh0BlYCjX3JJ+5WnHceDz6OKS7Zh3r3
ZdSHmi2tg/X5uY7AvWtDMP1/jzv2JkJMOnys/B+3tFBQm8mVuT5mRJXoRGIav994LA/MtERDu7bv
T6lDrIHqdCqghkBx+8F7l6tffCk2Abakd26HSgP3K5GyJLvsq6b0SdbqdrLPwdVl/I28RADCdzIM
n1K4aXAIXBjh4MPtF3IR2DeTp+NBqEPUIRg7j+hCxj7SuYXdSZdG/BHPvwUdsF5r7j2GeBLMYqG5
NqT/+AxRIjqyDl5IelGSWuytcetlBhtxFod6X7dT9FVeunv9yU8XwA4eJV5jqXcxs7kL21jf8Mt/
dLxZgJEDccL6O7wQMJhGN35v+dnLdaD/Z630xchwJ8l7JgApDtVnw5Yf5xfwU3pf7U7bq6Lnx92e
+VawkE9WLMOXpY+NROnToRaWXVcdgKzPWIjaTxT4F4PcCpBZZ6DKIffmc53PUA5VzDKWeachvX4I
vDbpivr3cy+kcBEzNiwpiOirG08UHEU5hoqGH2xDlOdJyif3DRPu444YKD1362J4kKwBv2KAGcqd
DoCo3DcJTlwhK1bh9Y4bOeLfxUeFbTQ43bOQjUIV1DKus0/OYpm470Ain/PdB6PcwOCTZ6ctR69J
VrDCcAx8nvCbrz3litfJfTjwA7JHnEiizfUFEXR9ZzSnS/D2y95i9oV3KMwSPadIUVneMbsQ3CiC
kyoDL5edOnN3VPoDrIOVnmb3oWejzrX+LkhWIsW3cwiCAn8Bl2t/DnkwAUk9S2FcmTcvbj57ferz
ASPlkUxt5C2JSJgJKjpcx+jVdGk0E+Vut8kz8NizNYg9fX5pKpXXZZPJo26gFcrsmtsSj085oAQj
Fbx5lQqrhY8Zh5fWDSxHD6a0hsD15D9tIIwVuplRANyY55WaRtBKxqqjCnJaMisOfB4w6mxsi6s7
61JyJi07lD2ruAfxqrVYlWVEGf79/rNd9G16NCk0a9iicncg7cgWdCIQKfk9rmUGRIZSzONlF4a+
P4+2HKqE2olJ3siHwh28PPV00V0qF12oVWiJ5gdOaLJNlRVmznzMWSiavQIl/xmxmE+nS5zU0EfY
jpGFD6SEkQo4nDzcx4nDX6Jq4eUmHeL0C2W0rCzrB8ZUkhLKmTJ68iquFD0GnzVh0PFrSeuOEpmu
ETWQiMNa+oqyUFRYOMwKdgtAlz3glSrKNrr7SDaGQfAap22cwGxaNFEa7kE3d6CqbTcP98HdMomq
/FMOUl+9Hut20l6w69GEj31D7NLqbQROypM6g3I44PVK2XEy3L7KxJgo4HqAdNJT9Ic+b3jPdHVV
/GUPOxYqLE6dzRhzW1YG7neS9mqdMTFcXoSu8lH0DuYkLJ12rqa2i3qj7YWMa6q9l9tNq4K7f22H
QIDoJPcC2kwsUyYvzplmj/n1NnAVpifrxnBSuSJo5KBPF5gyBa8+D0CpvhoBP3zBPDZtSUyQkNJ9
m6jWpgSLy+L96UShdtwPeonD1fQmS/339GI9qOFqYXOeAqE2bKe7zQJmYPOkFId150YXYUDsbgwF
hDgvQyD8Vn4ZWYp2+MTgQlA5ysThdeoDA6JORckzfR2ZlPZ4luFVc1HO80m7PW+aCM6bGeFMw8dH
a5yEXIFF1BPV0VNXaj5ojPpPVGiYE4/A4wf3Ie7SzA9gjtq2/nshJ3il6FjGshosy2qD6M9MeNxx
zp0YU/ffYx8rRTwJd9lFN489jYPcj8r15m9YH0DHcdu/n6M21sYykmKASrCAhFeek331zZz5GFen
zofiSfICWALKLnFOHMSfsua8FPTp/HUhlNLiRQsjqf45st0YsZrvFkK8oHmfX4tZq6z1T2fDC7K/
muJ7WNAJbYXW7YTHnwehafG5Mb2D4E7F3pikRDKivI0CiqmTnhTrwsskBaIdHCQA1Dxw8sR04qvY
I9bN31YlEHDMYXH7Tr48W/AkH7YnS2t7hVPVHH6mXr1tTZLQHquuXf+jxvH8I/5ymfZ2Tj0Znu8m
5NkVLmjDT9tK65USN0CQWRM1b9myrjzSZ9FS6r05EQSG1nbJGKy1oou9qBb0s8gQB/FWpM17FaQC
R5clA8ZvIsAKKDltQpxqVkFlyerkAT2oE00xbIzV6qPZxuVi/y8HhyeLCjNUth0xLYOA1XBBSHRT
3oQ+e51g18kfnEtG2+3rn9exHM+PJl+qJsagy2rg7RO42WM8Oy8JxLPLZjHi4ajfuRze2WQ4HifH
O+PTTdAbugBvgA0BbnB+eK+/VORxTw1l97aWmTve5X0uHUKedjMvfjFhlOn83q+gr5k7SfVL954+
TY1CaYgV1u6jUxfN06tAP6cbaYXpQDdmyWhSrl/2XfN624fzdWBb/oRj4mzs8dPg0Lsyy5ezquWq
vG3QeMW+wpkM53nN6xU0YQYOD9D2TtrPvAtNhDUNpiQFtsvsunpVSn3Mpu5c6Yfg6z6IOwe/gHHq
07KiKlzhOBb0p/9DMrHXqUx7yo4mbRUplVPek51Krl77+7cAJC8jkIgpJtzdQ981gOvK1PN4qzPi
KqAIbBl7wfkRzuF6uW5bHa3Sj1YANzCjgY34V5Bs9jzNsfAbSyKeWeq8VGH72SYrbk89p3SK5vz+
Cflc3zUleTy1AVDYIllpxMtSQhb6yq4OCtVTEwE9oLYUjADuBJKSSs1ZAlUqRR5991Ppoz5UsCyW
2YIB63YdBV9xjbR+3lHutE6N4LC1Lj4LnZhIbMqKnHMbgsnTVEOjDOuYOGuFRLDT2izAm50sn9B3
I4lWVM2XaN6luvMcsVC9z+hKxgDqDKMcnDZY86j3lu7cAAjIIGqtu1BuSvx96wVRgLL2t2sMIHXF
7O+PMANNzIULMG53tDVNjaq4mB3Az7VJRCTajBiQg4/VO8mI7m/BFAdBWSkE5RKsEd6F+aEfOgae
i79pImVqDuxhXWwbTwxZ9vNUe7N8PT9Xdle0k7W2SDMjfhA7tPbACT4GmESlxiS+D3hRPWCyyUpt
OHOwZBU/7BL5Y4dR6ikBYkcWxdEZBXkcJk719e29Uo45C0xueXYtg9F7sAGqdceQrR4WeESv4oY0
iaSO61GhfXOSVRV+lu0IbbDiWSUYIrw6t/MJZOtPwfMO5XsPyV7E1HHlhWHOseYyk3HFrsZ1nMQG
DyTobZ0NMUnNxtPxqAD/8IYgqepM1K8zQ/7eRLnjn8Lm/eK/kJ5y68oCCodLPNfree6RTcZDVjCM
4wTrQ0jj/7ITd11iVubS69P68MUAVvmjBRU5fXjnfo/CwLu3SjugPKxTwn8wlaQ/N81K63H02wDd
En7IJ6PmstEFclUO0yb6rS5bo+I9LFRAqj/VObnOiJEu5m0uDBj7JMtgZZ+3t5zNgznD6MN5TqIe
3DFzyQiwEJfS9vm9KJIo2MmeoXK5e3+4a8JRPnrRF79oAoGg6D7XBb+ZenT+6NWDkumBi/fChsFP
EToc+Cd+ELySK6hdosva+m5TMlUE7lW2MkIEm51aMujvkn+XBLtboNzYP6MN7pmwI2Eno6rFNits
1wK2TGEdEvbmMSZBuJ+ylOBFD4lNHeKN0NDfeC7WU6V9TpJ78nudAekk9293/4h02InGc9ZZh0sL
Uqbbesd+kV48CO/aPV2epEzBprGsoAlSgFvcV4uvsE1LcrT/oNPgeeWcazGctarw1ZWlm4e0JSb2
rDNu0yho79Q8n2WPF70e3XfRnh3cPdGmJxr0yZLND9m5jHylDTD9ZXKnC3Em0h0//d3kyc0yNI8q
cxir7HTaV/lNHI8w8kG1FdG/hWzdEVtTfCOp9If6nk6JqLhBSzzUIxfWpyy5v6lNtQNEk7lckjxr
v1X0tIWfzQc70pw2lNqk4LomSv1W/Yr+otLx6HlIzaHNnBDoZfbXlFoD7ReCzBQtP1cR45DjbWph
tRVsGyyrADzo3FIQ1tl1ugBYkwEqpXQZDdZri1nmL19HxJEjT8BE3HAKFgnyrQHxhQ8StL1uCcyD
BxyzssYG1fHvUCxeFDhZXNAuPcsbX9MsY7aWYh9PMOvlJWJ4tscIjojEJs/FlkFFvC103h7CRDZc
gkKYI2ZY+sWpn0FNDGQRKWX2AYIg7YOOy/yqTshndf1SWq7nqyGw2l6kfBVQCDrHdrsx8YW9swcr
ZuKMWRI0/yrG3Xdhr3dzbxrfsq7Tkuf94aXl0RWD9tnn/6NDxDN81lcejqr78SDXvFiJDsGqpwWY
I9Yd7Jbnf/3N2DIV87yeP33XkaE6G+GTjpIfnwbInslGp8OJVrS5NhSoL3n7/mPnU+EN204pnKqj
4vpnrJIbczeYCmXXiB4wcLjspQys952RYD/VMD0O40dx7j5s1JSzRi/ECqWN9lHaQQlCaNKykW5k
c8ZnErpTR46XyNKRLJdi73lx9w4ea+KoJUjv3J9m+5HSF7aFIhusk1Nok8aKuPSoJabz3nC3kcGb
bF+eS3LkgFubLdNszRmW5WpGYTlQJRXkCuV/RTFLCpXRu8NZ2Z/Pv/OocJUt0zrshEQHpLn9Rnw8
urc5o5mUWQSeGBLqX1Tg+5R0WOeC+XEXL6Nt4a0HpkoD4c2qiUjIkSIixVGH4sP4EevAQKXvz5w1
l3UCS5TLttFqPBy8NgIFeo8aB2yKcUyDpiC4EobDeU4ksy2mut6nJ5QoNX7cXW2zqfgI3VXTnh9P
0I3p+YM2sk4D89lwsDl1H/XNdgNmm2Q9EhXAMb51j5V8K+A/iL14TTprbMSuiNGOJ/IrBQ8gQnSX
Mp9NROHXlIj8bB0zrqP6y7zClMPsYIY7Q99G876UwsI+IMONKQmdUthmoRAhWOCYqQD3hX4Gjzzy
Pn55VhztaFch+4Aact8Iyx0nidMZGF1+pYIi4yR5B46I5Mx6RXxyMaDrlO2YXwPubtl31xDUdBM2
w1/OlIht0sOpvitoVIzxGidd/fXpWAhr8C6Sj4+9PEF8p5QJcuYJWKxS5cO/PJAxre4yjOwl5hMS
4s9UmCg27SQPHGLF+lC3Fn+E2RCik9RptQiPJ8eZ9e7rDzWTYz0MtV1LzYndY8TjI+CBG3YCxfyK
25jh4IuZVtavSfLDw88Nx/YZMWqe/TnGyZwb2vecs3aSuKo3D18hcLrdfYL2Npgw4wacf2+vY7/p
yFquL14VEgxUishHQpsBD2qv73bx42lp5FgAgHlljRfBuqAV+TCDU7va48eRmHq1E8Yi6rLTNk5K
gpbjvstamZwVd6hIldnLYtiEmpdK4i8wPH4nqy71Xbei7dvIhaJohOPibo8fLkR27i3Y05/9uqOQ
kIzwU+BzMqV5ToPUZYhDv7BiR7oUn/le4NGsiBWw2bbwv13pDzkRtoQegxiESl9TXHZsOjgZi07I
e8Za3sHeLHDUos5pbW3003vBn0hL22BpIJg8fhy6oPOU6xvjYZfou3hgNYV9hyAdqySMer5EU/gG
lr4c14sUg9KbNqXJuja46c3VTMMqPM32d55oU94eqPipESd4dXvMT+US/Ka57pWZMgSnuUGkFo+H
B2f3lccC4h+SpSZNkgWtcMy40PnPR/BoiOXC222+z95WyLQkFFRtBRAYUHGFzsXDNwKH/w26Phjg
vK9qxi4M63LnmvGGQCcFGDw5mj+pI8fxEWDb8WzB6bjVhb5ZH66Zrc7/3fJC9pjxSY3XOktJ9pJ/
raWQyArh8oT2GCI1Em4qfy57HAIxY1NQeIC2mE8+wPTKEDGgUYJksXqMrxTg3CoNhBH5Sskhgx/q
rmP9mf/1xb6vlbL95Bsq866l1z8HfLBZnFVT/WNubTgvYlyiY1Ql8n/TpYrATbhmOdkin7VWHAGS
FxFQboy/3WiLeA/lMg5iSAwBU0A5zU8/fO04pwcGDbdFrLDdrK/Q9HQb8ZnUXWOEGHUUcjFxpBNM
pKlvPNWK9Aw0cOII/pQqhDV2xijDDPHwuZvwJxfTGMR0/B78UNNjA2qlu/gQ3GLHdgP8UqjGSE4M
AY4XfnndENR9K4PNHW3iy10ZehJ019UmAzsbyS9kp4MOM7UyKvBtauV/eRu7fPiZy7wgctzZSc2/
UBEMaI9x8fEOJJ3GfuZdUzoiZCF/T6PyNtqcfYN2fylNSwvv1Ma9Clt4UnqETMksxLU4wThwZCke
LsCaKr7sVo1IK2KgpTXmZ7NY0hAYC4w+Fc6z4l2LO9JrEILI1HnkTCy1k1xispD6RgKh+xMSon8v
YeIc6WDr/2iYZud1cIbABuSEUnSO3LjWSP32s5XCX57nrnDNJDr3OTakbQ4vg7yWkK1fNtFBAFdL
fhsrbI2ybBrLHtYp+HtFSPFHf/DohToSadSb22q2w+LnP++hfuGtLJQQvrrPWZUcsnbtMakOvx/l
uUTyichOGScB1JsNQyZ3SVx9Uv3fsy57X16GtIke0A9mZ84AhGC16EsJvPdrYnGYeP6Hyp+wGA0o
U3VpnX3WOJQ6x9W021oDkF/6nA7T/CBqdPn+ypkDlV7eRXDWzU0QR5HfLcLbrLkpsuhv+AJ/v/7N
AlaHIqYrtgvgqu6Yzb57u/O2DP4kSFK9TEdplh6DNGi42MY1VRQi3PAaDbyEfcAr7otNnVrehqmL
5u/1FVsqr9eEeTJX9rpsmUEd12NOJGcEwxjcDJmYIGvOSHJOgeQ6G/+8oJeHAl0eRNMhV861tCxz
rW9tcR66/uhOqmlPeIBz12zIUhXWQJkIzfPcMW+3RwFN40uX/FdaM6foZ3WLCrXWSJ3JNAPZ5XHb
sR+jQ1QgdsQFKW0tUY1fvAPcF73Fi7ktKcdFvP0/pL41HcDB5o1sb1vxDWzCoa+8wUHjJ93OOmfO
DG+kf7qC9JPaIZ4hTMnFxv1FjS/NMGC3I6LENxUy4d6mV4lWRx4QRsk9VujsW/cdGcOaDAE6ZYeR
g/eAlW6PT54T0J+nRb3/lwqfs8u3pJ+E3BwS/kPswhWXfxjjnZdMAPe493+T1zx8NDqSpWWtG4RT
l8hlGyY78PEm+vEsrwEswkh0aUafL+/vJUxN2dcZUcSUdvnywQcUQZyf+8IIaP2oUhfjkxR03rqO
XXYUJ1Y0ERF7p6PRBZ+Q+R1HVcvTt8RAG8A7wPwwCLRi6gyUCmnvuGOd3mysseFTY4i3+OkJKxWX
SA6qV2oxvS0ycaeNXO1gvOI+oB5kDFVCESj7xpUdPB2tYetvIuOOoIjHrYKURXe70Ug6ndPidUzF
WgwmHb/1kxtMpNFc0ZeVexTI5uzD5D+2UijxYb2jJ4MuqTrhne9cXfX2axSGbDCpUU+RJHEezz/q
azhQtExsW+MVByf95tCuOU6phnXBrq4BkCxEfrRl5Vs1FhoETryEmvVgzimco/3lzMxZr5rKAjgP
ytEprEcM82q1Au6isV06dLVp022aq+UljwsmRoZX14Wt9Ps4fxgxf0UVpsA/i1vvUa2cr7c3RpGK
+MMVDRQdGjetzOwyJYVYHqDocyRKpbQJ6NKZP1OsWq6PL2kVSyeDDXN4pzWUPHo+hLrXmewNld6L
9AnmZEM2b3GLYFsQFvGsOPGPgyxWFKnXL2qmPx/l/tBvZHEyyr+ARK8h34HYn45M8SERJHCEKV9s
/aprBuymeFmmFWgNTH4y7oiXoi70TY1ZTSFXZIilF+b7Ce8/NQg9xmFDe/mS5HbmoNSYJ1wuuU7+
H4BObSCdWP6S/Uce2/pUv0pFxk4uXe2YzVGzYPfCLVeucT61SjH7WJMRm8OGMplr0dSFuM48ufZF
/Iefd7xQ06lsLQH6+91uKGFRVW+tUJD6JCX3SzpXarYjMqEr3E9JDqx1UuzQ/hqwoarSsqjTzn6b
b4w6jFpMU/tEwcw/kh0CPUkeGa/aSitBMv2hppqiwEs0NUsW1/XrWPK5S+G+cSTocIMigKjse9wg
XsZxvaxbM5nY22UdMqnZ1fx2xVl2qekVmPMQtT/3Jl8z26RttvPTmmMOrhd/2VexsUXDhJlcuFUm
cq4QiCr/nHXNNE9quOamg4wa3OXhK4mU/l2v4eo6qGKBuXVOmaLCtlTUGjwWPES6m/A0ST4e5ia8
Hs+C0OjKdijVZQybzyoSS+6SidlX34AX98JEefzXtbeExaAmCbCveQQ6bQFi0Kl3IP2Bz4hAgMgZ
7QGek8QPisGADwye+U4jNin+n/C3nuQz+4hbgh29msJbk4IYZb2ZABDIrWxU3e2m6coqLH2vGCVU
ynXef3kz0dM7ou3gXZyvj8E7Ux86wG6p7OaLRx3vHziGkOA4qjN8u3aMP+CmZhNqSSLYsPAlC7+q
hLuRYEgka9DZk/mJmG6FQkkjT7O+Icwy9lpXCBOQEpqeY48FQ5+bVOtMXdz7I58yxtm7X/A5Mseb
U0JuC6zk2cT7+W46nxZiSePs4oc2F4d4hu7JiCHa2Wnes9wBep622TMPw9trhi0N/huxEh+svA5Z
mrXAq86tWVOMh5MR6kKis11cPGBGCqJd0KF3srKnxKYAhx3wJBVO1ZCwzClHeiIMCsf9WnOJ5n3a
NfEXALhM0yPaFe2ylGEbJ9jGDOLhX9OBYnJwkIFkgBg61NiX2xYVPs+KGpZAKaPuRjWkqjspEem/
qMrhvkJtYWFIYohViuFxy5b5p7cGh8qEBic59iZFU95K7jNGhJYAhIL/K7TlVMHtNmSdaRiYvRak
PUFqlVoQlPJyhmsd8IOK5u2c415HrbmhDPCxMLYcD4Nd/cL26kPd6Grm/JN8OcMFk5C3JQ3oH2ET
/UobW3xQVEx/svASEXoEUwe3uHtZ3wAGQU3UnIVC9FuEpCT8gfTPXbWvkgGKw8uiCOtKH56gicDd
RNQ7lVxhxbWEMqbnC/Q8DHJTh4xmvV1xtxYdr96X0VnSSmfO4vvj0klh+b50rJOSl479ULw9Qgrf
aLn2CZuSlvnxLx457dFuXqcwfyzZgp1hTteA0J7A1eKuk7PWrW1Blt4uLMFhiFakVnUJvRlHGs42
vTG6ndu5x4XMxqfri5BnYQ/b/cYVIcfy/9D3gDaQ0kB5uQ0wCghBDKVjF/9QS0f9eQPdvuizjHwz
9Pb3OU9O10wyi2VaNewz63rtopxDdslZ8kENA6tYHQH2fXuN4sCCeqDlUScAuLhQMhjtAYYvF5X1
TqJHsneCCdn/hpLHh4PIZp3USxVdN83l1T60Bx/FL8W0gAbVWMRJ986RE5nA7SwBXA8JiBefI8KJ
Vihy+W+ArqkVQ4wGrFOE115oQdmeeI+53b7GOLjAldKQnD2zFnzpr9i7CN9LMdSRgE34+up1d3ds
l2Ea1+WF82b/nUoGOuuMWTl01bdCRWfzO/urqNufr8ea3ihuclip7fsRjzSsoOuy3PqioypISxOn
+S46z2gX0GopXd/ntfq1wmTAmbQ+JLWexNrxRVoL4RLydAjBqlYukrny67RAntO3pja5Eo+jeXYg
AF+mUZzxPTNXiW2UyX8JX/XQxnEd41uj57gPJXWtdAxDtM+Lbdn4a60rYTfHXsRrTgiBZqEMA8Vs
3EmHDbXzfJWUlBh4hXDskOXsIKH35FC3IP2M8B/wFzmHNfq8C4hiyc4i9LSqfcdtTTndz0DjeZc8
29ZXtiuKmutvljBN2Y1V/GzrZxG2CBg59ieTcKeD/LzTSBw/GGUlPCDVj5eZb2fiWZemaCk2vyVt
2p57k3kI8oMahM7PfF0HNjXneZOK6euUUB8oUAddAPvmZqMTs70pSuNDoLQrvYibTq+rc3ruZTZV
ztLvXTjJqzi4/Qhw8tRUxxpI2D36SVMXxqsEjzppSXdSeWtO7wca2yvqq8grkgVQctrk86sz+3G/
4WlRuf8RSo8Ia3kkbbYk8ECPgdBaGQfp0zf6PlFZ8AqS9uqLbCkxocHMwm+2xdXbByfPKwmh49LV
xnCuM8LOo3XK3cqd/VprWKnHE8cO/VSv6vjBC0JcuEupcgTtvkmfr8UVlkFlqZYRBwBdfbo7Kja+
Sfw7VLGFzAemuSLAjFhH/Nm4spxmiDek9iCVF/Dd9vB6woywq6yJ+aWdrVQa1yGUGwVa7trIjFlF
j0jRduvubFKpxrV1E855FIUtAXq7/CSODnSFtSZsup+4z2/oOIpXYcucOST8VoTDyI0SR2dAL2Wi
jSxNl0WpOF3KSYm37LHR8b43xI9Stn5oFflTy8bGVbrHJnAEZppqGydXhUO7CHtiDHmiBI8hJnBc
lsXuSIxVgU8Xg6lLC5aYpfj1ykX/nG+jGe+CCXIyblE/ZqfoUKc2w+H1TF4iChb1Q3EFuII4Ozzf
Ztth/F97N0hPKxTjpjpQ1RhsE0odbO3JMcazuM64HrcmqrlphXkARzAKLqPRzdKt3EJoMFYKOonx
HauYhQwtthZlH71eLGHnENS1eshSFaYrGrBUqch6qdThcR8L4GbWIlo3OwHhhDXPc5VVh6uuhqMl
6wnHUoJSBGvRdXzL5vOt0ZOEYFvLImJyH9X0q3D85RmEGvZSH5lWIAQLjEzqnjypl4oFIDpgJbcl
xQK1xN+Okxi5anLd+ijvPPAwS1laGOUPN23Q3HnVKGAzZMJf54qniqpUnbHQRSuqBhZgd7Z5VyC8
XsjrnYlEgdwnKwMgbCjVQ/ekwlm1gvrXYnGUyXZH47CkvUE1davcYCpRewVhS6GC788HT4kml7FR
slg7q4UM3q234Pq4rV/85pKJcyx31nwjww4TyfGuE3CYYK8Y2Qk1867mPg635CPln+wCLQHBtF2y
X33muofgnbXocwMZWeGSVo5FT7QKu7mxujs0Xg7AEqpsifPnMqkcmqbXGSQP3UvL1aFmzEfw54ac
MtpowlH30b9nzrjtgk7B/W16dHSJQDomEUT46ojr0fY7qCxLfHhjJX+wuaYazBIbBmtcRgIjSYSM
GeSk+XGrbt9jyL2RyQvHMwPDYrSByfzF7k74yOnNGR6VkZjo+vT//DwH2/6NzWElmXJI61CbyeMx
poKAkvQenEP2s7gLS50twjL1OODGQ7n04HscO3jU5mTecCGH11rXXtoC2pUXrxuYqh8lw0G1H+xK
9Kp6h4CjPYjhOq1i6ILTaxN0815oXwmnaiNFfeBK1rh4wXl/nUhzi6DW3k4yovQelPWk0hTJ7A2d
nJizXx6AyRAPotr2PJXK+c+jRTAg9XfjAOMsnnhveifRMxKAXUbALoUA2eaDbtWz7tjDhrL5EJTR
m95919+2n6Gfhy+souQykrDm7Rwf9H4SOrYSB13RNlF7Ad45X06ei7D5srKZjIWsoT5fJDccU7H6
p3VUoAE3iA2SDngpPo4M8chLIFXzA9fwDZCawCzN4kH0b5LTJkt3Okg53pfqQv+Dg0ao2Fmt948S
ht+a6gSEQHuNWCfMoLlQY68yzDCeJRCJFXfCyIEsRd9JccMQmJwz9s+22oTk2wk3f8NZX3CiQBwE
2BEiCz9568QQOp+lI0YrMspeGnIwfiiI0rR07DP9p3WRiscCpmu+0wOY07Rm6jJ2IOMVvP+H0gEm
3faldsSBs4liUzbKrF+BkRVI8tOjS+HEaUWMrGcXAp28bLDh5r9k+311LbozdOdcZy7B9FKars7X
3VhnQMBdwbX0H4+GUNx9DL2TeJ3XzN3QFMJrn+JTq8RwSSuMU2xm+ee/1Pa83lvA0LC49uEs3fTS
p58CQsVZdEkkMosSeeHwsxkvEztUfOZb3wUqLsNvDGAYNs4loXaFFSf1wfAP1OrFzh2EBX5WeZEY
pkr3x9DwVNKJa3Q0Turx6JrT7e84Pp9aVa8dF4B0vkaz8durQgyDaDWPZywW2MfsWQgbVyJC/p0u
zknR4yT0u7SnKNYSxxudz2G1rLzttZdhg2ZLo+ahsZFPl0U+A5jjTLXEs5EjMJ13JSASdNyDtDvq
vGdtPJoH9/KM+4TnUbIkZg2hO40iKl1ujKZbQlvXF99lsTwdWBmraffAsMuKps1Urci8ITpYha0Y
DzgxSVMmAQHRMavYgNAv+wS6ynuYqkf5BMJapUKc0tMbQKn1TfypibcFHwP1ZBdVrUpLcEdmxAOc
yoTcNuJDfW6lOjPy8TlqRzjJMHQBqnxbT5h+IfGLBYbh+ODxfRgIX6rTOvn5uP/egZCUC70Aarhl
2rOxRIPOiFonK5P+3gsotpYnK6dp6akgjYQG8rHqxm34ptzpgqW5HZGerYDP7sBpk+i7hYA4QCld
+AZu3i2mWAjtywsjPtTTRXB8ePfUlJpErHAYjJiK0TDn4HA5ozKu65uAUjRYgpdzsy7pMcVOt4hO
ApjXRSZagORQ+UheI099ZsWgE3JxnZq+/m8xDaVoheTJY60VE78ADxA7qtg5TB5fN5CjXfmk4dgb
XQ1DbKr1xTgb82egLBG13WtYAmbeBRlCXaesnwgMNHFN49dHxbeYZ37W9froa6NNrUN41sdC9F4d
PK0TaR6JzwdMqkqAuIhrD4j61cfefNOqfVtDNxjRYfvsSJiwUjSsK6MHjC8GtCrY3gkKl4V8ZoJu
rbVyO5rvazfuWVKUPOWJ8uL+GpOPzIWL43Dv4E/kSH2t+/KpidrPtssRHGYOQPCCzyKdF6dFoCln
hnuQk6/CjS9JnBQo4wzaFiyf+0eQ7+PXzbD5cJTESf06AnxAWfVQE4lDu3vRiEgsylhjLM2+Jxvl
lLWyA3xSYk+to6pqR9wnBAT75hKQvtesSecss2STIh2uV8epzEmRvHKv28EzLNPUxt+4vsXCrjWZ
E8jreCl3PIL0tssP41xn97l4BiBXuic4VLYMq5QyBvU4WnU0TsFvL1h54m63+ivb3Q5F5t0hwXDK
nuH/g1Z7GTHAdqGHpQE7Dsp6fQA6o4YsW1DHEVZgTsEPS8ACrzCoF5vh+bT9fH03h83akEf+nuHQ
MS62C6rBIU8Q35S4KGCjzCxiViCYzSY2Ucgn3QFCscTBpA5P56xtAQOVDsPlrqgtw/V2a5WWWrq4
zfbKy5Gdue5wHgDEXI3a5nF19CXFdzAkVieP0/Vl4foh9nub/D5zIJB8wV9OLc3Dp6rhn2LIwR6u
ZRSD1qGkevirhR3FKht/qpcCVDn1d8iwG1mGn90kA3TfrDhfxpBX47uVcr2T6PMG2tuk15wHzMfA
VNRdIgyJ81FoU0rnIapDfCUTjSPYdBj/pOjPCHQ3EE9huZZWyHZHoz72Nojksx6rR00/iDZJzeX+
oV51zCgyAS5K+IvS0wnjIwM5J8tfEsn6CeiTRkXTqCloDnPArPjhSSh5vrnRx8mH6qXPLTYeTYkR
ux047YOOmf2tflsorq+/paT5gYiHqKmhDHidBxyVabqLMUCE3dSxOasgLtz43nUFuMyluQtBNY9u
Dj1SC2jXDmRKZnMRuSMSSTtjL8dYPEA777WMHNUvePa/+hKsz9LG7nr1srHj3AtJzliy7pGLpnPp
+Ep/tXmJrSy0T2wC0gKvlr5IKWpNzzK+PjTz+cQPznEjj47JGE/Auvz2cShyGjWBpovsGCNu4FGv
1RyjlJ305NgxARJKSifHuvuRSg4uCrDBQ3nhuHRXznfF6fYGFGVyZ0NihGZMe6C5rVNg47Fbsf3U
cCJ3dcjpnG62oRAWlprMADpZtUd91sh8l/GFDMUZeJJzRBry/DVhLZHu7njcHhHIaaiIfeUk7cNY
srNyH7WcceI0VpexOjEtM8wtUfPPrTiiqflULxhnGHgNv+76GNvHIQvDCQ+C/q32+KEfl/IBXoCo
jZopwTSVKiolGhA/gCuwpzVNHVXdm1Anh/PTTm8XHhKmkxhyZBI2hW27PvnOXB4mstjmC+OsIW3F
juM2Di2s4BzgdyNvlp02cp+ZjpNHnj3sX43u3/plYJHiTHmkGhaFFqI+V1LRkCNGTDlzy7qfN7cI
+Lq3xCYNJKFJkqn+eLM9tVrd6fefrPdSWpNEmbSLU6tXo3mPk6zFlhRWkkk+SPHc5ErFUuTZw21/
4Blw1P9l0H+HdUvONWajtIDos05UzJocJBUrJFgPlNAfb08zuT3PLnnWfuXDLFeSH91kGjPil55r
barBuI4HBpD6vJaMNlkxA45NBxbUSsv17YAUV/epxfR4G//gLwRiqBFsuCu4d3uv+9n4kSkoVFMV
R9biQdxjsVwMk4rVnaRO0W31NyVPqwnbHgf9rxfr5bgHbmPqB6xOPYSUb/wki6L3potCoim2ld7Q
Eq5PrpmOPUedNNKrIqx+Wj171/tf7OG/U1GPHuJb+9x4GnJkOCmvfGlj2ZsBeqFgrqbY5bN0v4x0
+sEOOz/Fhz7f8gBSpXbp+bPhLba3jnna4jPwZz4JO+JhPX1DOP3s9XF3UUeKC4aAHdnM/jf0KqYK
jBY9c6Z7nvijb6zH9cyTOp8xoZQhxyFlFpWMvZi74DUT4k9aTEvarerlu0ASJ41u+FzgubnmpfO+
+c28iPdHzw0kv/e6quAzpAwU4St6cDjGyLfKrqcGB4KzIVKilcFscOsQ0DGlwIGSbz9Fdk7cVPNW
ta7w8xTO0+3/TQygslhcBMzhqsZHzrNUMAsKXdqu7HPaMnN5NUtx0vFBT5V6btoXUeSHeHI0noxW
2oH7ter4GDtRZXaqLP+j0jv+iuwIyoGHAVwfQ3DERZPkIX+i5Dzf2jlq2dtVN7yFGYMLw6+KTFFM
VpAW9OaWL4JD1DdkfVbT0uoILI5UitSIxIQRzIqZJYtgpcM24Oll8kxcrm/Uw2+GGj7M51bGEGl1
DDlLP4W9kCYwjYb3zmHupW/BWvkkyRTHQ4APVwdNwSB530arPbAdRNXgV5iG7feWi1UHiP/e6lW5
pdD8l0C9ctJmq4FlqZ2JlGbV+80ht/997actx6mUintWM+9ke6yI1Bnjd5YvaZrKu0SiRIobriuT
f5Pr4Ql105/ndoH27mOLr7hjIq+OAJK5yluJ3fqDO18jSd3/KgEEfeJjvZHDfXggjblN/K2YX/wc
GUIJbDotFsfmwnfSxaLXzjhHxlsepT/w4NcTcxuKIE5/Rv5bux7zSx1F8/q7y3Umf8Y13s+yhZEW
DsNI7XFFMcPJFmN/i1X6Eraadmpk+bqKznc/KTdjebPRUgOd0u/Vl/eiFo9xAn+5cagaa4eZn5EB
xfQ2kVx4cJzYAzo76jtrogntgoh+AlKaJOJakW3MF99KSKMTRxVye0U7N+ItymviS1oSyq8J0eF7
gv6LKJa/I1FI3XseEKn8NYEFjK6oYw4+7GX3Jc6NdY9PYrQNCBS09PYjw7dEQYpP/NC1XDkev/Xy
1fLHWByPqYIxFN9JlPcctfkUMA8aAlKGDUqt/OLZtJ8EcfoO0HjJefVPU/iMX5o3nplLQm14apDr
P2ORz8U4BwzuypVKrUi2A5eGwkops7EAFiKuwROlSUPifvbrXLteiA9tWV7FlCKj4qQ7JZlrGrg/
zMB54WUSN/waF8aQNEczUeeJmdMC55daw94Xgotia8Y6RGcJhVkfpw+c450gsHh5iWTgkNkW4hdj
C/yRqIXv3lxsLMN7+DEsTH95ZmjklUkpq3JMHOZZGAH8HukgHIl0LJeOkpBnkF3fiTjMUnjAFHHH
gRFDdHLOKSGUewEI3UncLrX7KB9E6YV3bU77A+jkmWUKKtnWedwClMPKlMoAi7RM4o+ZjWZLzqg3
YdWbS++UutjCEW/WUHbuSiVp3ATSq/mMhEBnFn0JqSHsR9flGQfy6oypqjaBmrFupxiKPPZeInWS
zYE2EquriCuBtV3i13gS2TVP4QOvjW4X5dSGCApwTKXX5XpsjcXv3bwIdCVNPE2INZxGzem9cCkF
sJmr0FGPSlH9kXP5g85qiSkC9mOxsJyo4q5sgrxuNsw37S9Pi+o5x5SIxliqCzoZPGybCRJTeIQx
KJlJ4XJVQl8CXX19+2o4foqpLvQSRJYfm2AK1G5fVXPg85RhnBS5Rj/el1MpSSaNgHPYnSS3B8HW
CXyqkiOkNVEhL1KyO+7m3OKD5PGmzbA/Xx4rjy3e85lMxyGkdWzsBXPB3HWHE66/cp33FGO3kyyp
AUmM5wlUw0oSGTKudqvRhk9Mhxt0AZTW471m4TTSxJCkSf3/Ys5d5icITUE+hyV1fsgf67aicC0x
u7KjJgBxuOGSSz2vHH91MCgowjIC4OwtRy/rg79DsSIZU6dW6dWKOyt5mRsEU1Dqb+n8+l34ZpfI
S2KcOpimwML0SeZtKnjasreSi4WrlZbWjF+Abm7H1WRp3nUr7ehEGpvWxkHrUUHhtKVnXJIEcDxv
rrU1aQFxJbrKiLOKA4r/l8ktlKp28UCcGPpRnPQd/pKO9mTWFxU6LO+z/K+WfBT4MFTIRDZgy8Y1
XdZfLIg1jsuu6SJjbR8CGRILFlCP35x/sQaqFbdHBNn08arar9YZch8T2gHqe/TxCLgpUpNiZF5H
Eg4EAd/548L0H2PXHBR0tuQPqv8RBWjMkLQgqre36lWsJCFzut/E/2zlnVJmlcuY+vmm8U2NIjXf
djNCSgFTmL3UKl1MVIpzTDwcbG4LX7BOPjZ0pfHcCM2GvWybtk39+on3UoLS4Evqa7Pbo47J34Hj
JK/r/be8OccrNFE1wIRhTpBezLWFBIGolFxhw1pV5YhLEsQjBbVDJdCVe4mbyQ/TgQZxteIfIaRL
Cm1i1zGsRYQL1anS5FPRLxRxxL4z3YKPSPMel0ptl9ab2yKbd/Zq101mNKK3bzwtNNeDCAk5G+bI
97z1oSRHCW1lnMbZsIcvFixT9vZmYR97SLrS2TNS0Aqp05bkC0p8xiYe9sHpzbudgJzd/b/AshXM
jRUwyEpH3Gk0Ye/sb74IeXOGILlBSyVgK/SOLG0+zb2Iy0gvO0kc8X6n2fLTupmS9vd0m4sEjdjq
vpceAPlBbexr6pGVv5Q5wjFjzHPguAq5/nKn5Xl7tq2JmHKVxGuW0a6C3RsyyOsN3eGseflAb4xL
vyRYgLoot43hZ0HemW2dZQ1i+P5P45f5iBsvVpwJxCMOp81f3w6SlwS8W/xaexB7QPSv9mtN1hxx
03pG54DX7R6FnHoTXkItGIv5ZSnrvh/G3k3sT4SyGz10P3+xMb0Prku5RZqCvXeUuxOE864Ow7eE
B7OkYXsMfs4qwH61XpcioVP6mg+SOChIWVYvkQiR3TajePdlZq7mtPyfG9PP9C8RiBjAdi8gZDuc
eg8oktDWzldCvfSqWcNLWE0kqMDnujC/P204MFv5SJgB7WU8P+ptnO13LAhDwm/04GJsvY8VK46a
l8eYMQKFVl11b4EjqzTGurTad5/sITQ4KD9AuSzhXXNZ1dVH7wZw8Uvji/bjc86s7gqw9hWeVKFY
t1I7E99zpRl0Fij4U+qjs4TAEtJLGDMxEv/dF53S7QvjtMvnntEuNHWonpydnMRCubbHBj7KtmH3
dodv9ojgQAmQpA/OwD2UsSdGukGdffdXFlaOzEiccPbXdw3aoqa7SCaqavQv1h7zE+jdTgTe8tn0
4LJMzSa4gRg8PgqyrZ+ya5rEeRjqoFpAU0+x9DfyPpTyZNg8XXfOIM2vR1LDK7LVb8SVUOJja+oh
E53XXyJl0TOMli1aqOzN9qmsstJQVhIK3X6Stpl3fteXXyVoG4Y3+Uz9JMmlQEiZ6K8ird0DcI3m
pqOIEOsdRCs5SunjmrHqL3yyBNMJdXgyxd37EQNHTdL21DR0JHnB2slE1ciDAENrgsAhlPuu3ysM
Bfv13V+84uQjqbdQyVsacka5Vv88LB0PUOonJ05K0ZlhX8L1gi7b5b8PG7XHylPF3mgup0U5jCWm
adCXIpwSPd1syD+qUeNNCmLPrv1pc72snoKd+JEY0X+6EALOctuBz6jBH8yoFE1IXwLZxVNxwHHp
SOBWIzf09HDYVsVppU60vCV3RCYTKlEcqzG08vjkhReMfMuffKOQFh47uMpHOqNh8nC6pPBIA7V6
wJB9X2BOa87ay/u9M7Y7bMNeOD3G2mtglUCZelESd0oEnlw4Q0vRU3uXwAClTHna57IsGNGngBBi
7+ZHeutjU775nVO/rjyZQ2uNDb2jyFKwn04CzPjKnNzQjN2S89YgvJAHJ6ao+pG066JB8VIe0nNZ
SnMgj3IOnKLHFBUl6HP61r+ZioiMvOQzPx5YxOwVwbuZremF5SE9Sezf+f+f/vSwg5lkg4Obgeva
Y6aumDagJfYdmEArbNrsgJzENn4NZEDh4N66b/ONyDfBrlsubPpQkDoP09YDrgMgI2MSYQtqRoou
/reB8nPEgI19ctcChH60UVLNcKBO6e4RfuRgb3Qc8jUqyqbfBpd3y9D8qDMjfKrPl6Qwk154cVBs
gDqOP00ypnS9kepSld7OTFO9D6QGLxSLlX4iWGb+qFcfJUw8ieSRFvuIlPG/5vSoNPXESLR6MqDA
mQ9BR9S4jalCsY/hAbSDzIkIRdkOmGmP9vuEmpvUpSSOrjPeK1jII5GZDMonY6GK4nMXK3w/PIop
33aM+0anuNR99ZWGmJLqY0njyq0Ms9jXmyIK40zGLUDFG/f9/KANyvyg7pK+vUdhQ/+E21H0xS0w
0cDgT2HgTFAa3wTEByRdFC+KxighcMBnUIfEp+15Mx8k8rlt1J/x2WIHhnXusmQ4j26hTd+m0TV2
JsUMs64rActRL7xYe6bByqKVRmUVYZqwq7RzuIgOtmYO4zOLN3rUXd7xBwTxLCeqRm3Ar9o2rVBf
QlXFRIzRqr2d9rKrVMOVQ5kQdSHmeLPZdeB30sYiWDIEyW7l+ldD3GP0lDwAToYHqD1M4puGI7mC
f4Ot3Goqb43sVUc8y0/EoR//yeMYLTlugycjYJ5SjBArzeWIu+Us8jrB7ufT5nkFjCTR5sfchjCa
Uctd9gIgh230dl8TyMqiSfabga4Gu2iEGdtRet0+mbhqJgxN8oDjgHEvRDnSqT+MHKhuBL6Tofdw
eDINs5xQ3xzVrST5S2X9V04J3G3zmvyHdJPo6zIHh9ygGs09+Iap/kx62YZcqqQyCNFW00nXJ5ZP
kokuo6VstuOOEx9n5H0oI1GAPaQB72IbEDJmmQ1uiaVwiLtWeSACt7GgI2NR2y3plrJHGYSu27k7
el39l5ojJj1iKEuvxkGA
`protect end_protected
